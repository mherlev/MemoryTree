// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:53 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
TQHPJYJQGRrS12YG13tmm3+jOY7XFawyRNtBOABfSAvhBWQkNZWZAAgWzWRaUTCz
vUZTKIppT7F6qaNx9QHyEXFwASnec8VeC7LNMi6Y7rrdpt48Mn0Fs5YKrSQQ1lqA
EXmlXoxJMjleTzysTHNSwrvQ6jVIIF3xltg7Slw+3I0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5056)
VJQhhL1DU5V9d7tHYoiQJ0sDNFOREmVRUdp7ryeO7JxDi7JRun6Q2BZ1WRiifwLr
t9R47eMIMjnUEoXiQBJl5yA1+kwBTYaow3ZxCA9HM5iSRmT8/iEhT2Km+9eRumuO
5o7CSzanZxSMRIN+CgjU7dHKWiu3OtF51eSSX4cc+ki2KL2hdVO/N8wHMkqrih3L
IW6ul3REzBn8BLo+wNsJ7DsA5LBmZopVrQhJS1wlZt4WTqEex4M2zpNViYTF3IVE
uEFXYr3b4d40Q3efqF1AUIBWg1Hm733iCUJX5KhcMZDS182OuIVLphlom9UAHY2W
6vztUu97cTuuEep69DarigNuxoGrpW0/gqevu1xtOEzVxjJQoSvPJpADeID84Ntm
j6ABZd4K3TvnwVRbhZ9uUBaZ3CRCWRRXHC+qHa0bt+QMPYPEdT9qIZBPCBeCXfaQ
ndgQ56Ds/zkM8SyQKqAOmSNxH3AwCQX5Xm2XAdybLmRK4WvdcsuVaR4nPQ96cp76
Kc69N6tWDYeWQ4LGfUsQISTsCTAeoGpWhcSUy4LVQ2ZKOvRtZipCG+RUaRTLXsCk
7ajEmBzutStlBjabPXA/+iQ+Tr2o+9Dl+2D3QEk+AbO0IRPh8V44SEh9SpBKrgbx
OE/Y0iHrhoXPxAMW3ebOO1LUjVKgD1bbrpPIoCca7SrV3h+2SF8eeV+dLyatuoWv
0rHP4HxY/RWVr/woc1eg/rq9VkIRn50nw7nmqbuz0y9C+OLF7HVCjf8m7MPL0f5C
kEgJMBm0mV0J9Vxtg4FB6M7WeGp88tWYrQZvJ63mA0dHiL3nP7p53/HeX4WBk/hl
hCZJrXEGQtIdQEFRUTc2L3QDrK7QbloSvGUkrbTFve6D5J0jyHUdYYg4w6LyXEfL
K8vQS5p/2Gs/gTMSXo0MWuNVTR/4sKlUt4xh53jaP+Ai9v1JXaRWlf2phmLpndX6
cN1Urzb2aGKbGX7B0Wsr0l2cUrlBpmgytK8bi5WRYbNb98m/9egsTHJvOY2Lvy1p
bck9ktVDYfUsNMMjeRrd2q4sSdd46PTYyJM30DHd1ytzCEaqaE0efgabbgJcA1Gg
LqrbFMTL/Hs074mILuaqKKet8GgLEtQTOl5sZbFrrZ91Ny7DTpc3ehRDXPxevn0d
pH//Zh9MW84Iyaeydnirr36t8Q+ISznu5K/SXzqXpQ3YzZG+bIrx3LZxXzcNZvyj
hkWeM3teDXfYB0PNf0+4wsKQ0fQPrz0OMGM6oPncuSz01G70FqUA9hm+0DKBnvzQ
6bIGgxUgx0kdD9eqgEQMxP7l9piZ76d4DNt6ngFJYHjw8x00wES1R+/OZo6iPqdh
2C5sM0Ngg3gBXVi004hRq/4cOwbDKfiPAtR1iEaOfCN0qUwxM3lGnOWqDrFUzSE8
cfy+qGvcomzkUOxbEkJ6S1iwFL3CVASzWmq8ilDQY9Xa4ENKopZHdUMLCXDNrdfL
F5nRHzlnoZuDmSasAPB/MnZCNWAUbl6hK6UhPcmzurSAgM5jWq+HvS/m9AXr/0NX
RN3AgWd2ArnJBztVnXGbRYtj4QT3GTkr5ZkhByvSr1P4Tseakp0MvG1Jxqj55oJr
vm0e1tcGBuBtMNpFjNj0kfI/v6xeq7QjqktkqEPYiSxX127kdfIzeqRU1IocXrgq
12nMygXCWePxGt2aK8+2uiTs1AbBCMNIin4JdwuZz5tk+8Vk/9fO83zek+QhJ87L
h9lQvBaORsI5xgYIUJrA560g921SUimedaecbtvkanPSWdftrg63mNFsHFbxqmnA
AhEaLJwZxtmHwBCG62oaC5MY425Xom8a1ZJ/4MMsHBT1xX4qLELIX8ZNqAhFCAHH
WXc6NqhHDfHFbQpg3354RkVfX6Fr3unw3/1Xw0QVj9Tv6Nz38w4NHLFNvhCesKk3
/ngWzUMAwDUOJ82GRODr8bd6PR2wDbmf5u04fxfV0hDEHonOr4OqPlVpDCd7T1nt
dZ7WW9ljuP/zxQpqqGs2j20L1qjB4roXUC0WpWWhigdrOqVaueuZ5EgNcfPeB5Z7
UjPPJDOmkW4ONg3uyFnbmaOZoma6iI6JSdAGUuf32lJvDBdaehG2eDtQAJM+7KCs
oGapJDur68t88vytSzB3DE9DZVIwl6SfN5titrHAiSeWcc9fprbwLx7fjd0jD4oP
ff0eyz/tugJK4sHIDz2p0Ev2pPp5cjakv4+xbQZTmSmggHTq4zSQD/3Gr5gKPmNb
VgbuNOw5T0MNY4tjlTyb/raj6C7sFWlrNB1v8OtZg3UFLloDVt0fdrxMoT09pAcP
3zamtsK2pceJQeuGCd2VSfrQ1z8Eb48V4GZcOy2n3GL1ykpTrV+ebjH0TBs31fgG
bGe2u2Tg3W2250hU9RPF9/3+KY3EFFN1TkUUBTxz7MRPjCArCqGHb9XLLpdeKj6L
at/vKIwo6e3Qx9/7IVsIWagV848EM1WBRXOLWK0K2WOQTj97V1+osnR/oJRlTD7n
WSzuzFNhVdgMdo9Ll8BkRX81ePz69KOx8pxL/KfHzK7wh3Oj1VDN71WwGQjpNidc
Y2XsdVRzmQ314pFVaQi7u9Td15G7t8U34d/dk42fc9NJeku/mmXni+se27d7O/tW
z7j7RxC2MGGofco9s7FUtdd69zkSpRYEw9zSq3iapET4OtKGJr98i4USMSiS8S8z
a/cqOIvrkcvQimUJrTZqlgQQYsitoV9vS00ADZrSLVUiPG2wIb9GcTRhH4fZRA6y
ZEHv4ELR2VBdOBCpU2AgvrFDX0oIOigwtmLHPJccGBAYPWzVoFy5a7W8CydpXevX
CtvLqwRcYBNvUEWaTip/JL8bTYVa9ZHxPGzRrhtyHcY/AuGuEFsIJv4mtYQQpeoC
sSicd52cG6RZTMY/8GsYg/DfdODLWUjhoaXLQhmAXd9c3bTRR0ocVyzIhyXTKRTh
hjjctSmObrELU3K26TslyRvLTVdbv/AkyfhGqrmsaH350E91ns8N+4d4rOslQeb6
EOJiIyVu4BI5HdjXXrImi8E9j2IzGNwFXVea+2FCMPgTsSgHjOI+D1sO+n26nY9N
/mObR1HvJA6IOf/9r7jgopsvnkqzorNKQPpWFphP0W3vUhtIh0WoABCtz0wqwLBC
tPdLMr1Z9+C4fInMNHmXxeCv9l+HQ0NQtPl7joQl+tuMfsVTxgqFJaTSZOrCVxs8
a9qOeNYGW8VX3y8GIFn5dWSt8ATZ68Jtf9G1cdsvaKpTNfdDE9Uec9VdcDS7z9su
YUg2LTkXv+75vUlwWYA1o8xSBYSjvvSup8cV9R9DW+N2Mq+oqWfNtPwm0IMViaPc
WWBI1em5ReYQyjdG0UOeyV+AWnent4CsGUoFUmXFWJRy1j9C+XrBFA3dEoA9YLUC
4+tigwFNfR9Y+cW8s88PvYGJKlI30zjTll/FMCmZUJ1y2/1kHl/Q5vZ50BMxrj0Z
f86jmBVYnitFpbS8TpF7znR4kiidGMWZzISwq5GA3JREzyE110wnvSDbEbA0FXfu
mESBoQBsdbwcEWzz/BoxqxRkZ7nWzEuzqtsMDrukx7eYRmNx3r7gvNu3VdTppK/M
dRh2FVZfSDhn2YLlzucnRMkJzk/WdWUMWGdAYe8o/xicrmIUWp1yOUJAO+kznrlJ
6TKVvjv9EQ1ZJHNrnaPs+Ak+oDzjQNLK7MeRZ9WOAct0qg6O+dqi77nsLu3I8R0v
bbhxEkkSpOCreDS4OqNN1Qg+dAVh8j4725jxBpOxvJ7pzzNulbtm6AHwyxyv5Gij
IFTvIsHcbAQSQ8+AKxdCBGnJVnqgyJ1u/xXH9+q6NiXbyABcKtUYGp6nf1Y+vM4z
XYmYY55roGyX5ExzQF8pdhOpJnVYxG5urC9LSdrZRivuIFwLnDscwWdRkKyrUNC1
8mTsSKtdRXy64ik7i8eMoGjwb1Ubbh1Ws8dBRGfhyLi67b52AMaHRN1LPHdLm9ig
dS27VBbowtoqadZ9Q3YJ3mvJ49oa/ID0rdSctnL2JLsQv7bxKqpIA1GsWRYHTVrd
eu3MA1fpmGbljhC01EtPBCbmSV+KsQaup1S65y3LAwumhW0L8N6AO1fuoQvwP93S
9CwhoJOfJcUwxIgWw5PonVOgMXd8M0dWP1XKClRp2k+RPvg6jbhF2wOVeoxRKnG1
9n+msyRwucxErlw9GGhLHPUTY8iWzvAgd5dKSYGpYWKEcZ8234GfBUk031GOL8uO
eGXFkaxF3izS/WcOOIHxhE5LW9QOv3xWDNcZtnIoQuLdlpGWGVli2o1EShgaVR+V
u/liOf9HaNM4U1XLS/oSL2ad0hpSzB+DbwspD7g0FonHzygfXGeZUSHIInszMudn
ytQUCsYwuzEQ/Z8dlPVq6uR/CIGK0jNeViXf8wl1sQJRFiI5jHJjl2VUMDYZrcXp
f9XHuNKNiCVEip3s91eqIQ3XmqBozdX7Uk/GOTnNSmoVWp0+flx0cYRyiarmVWdp
IRMKtwxem7T7gxNwX9bidy6NAEmc9opCs7B8i28hDMZHWaoalBBg4Vw7qBLrUc+I
16YFiFjMGKmm+zuggm5aDlvZdnDDbVMYEgEC3gIzqQ/k9xDloVLpfkQkq1zQdMYv
c9wqEECVg7bYMGfCADdCWySG21xNGJcR7f0OrKCU3FlPRDgoTmk0ZosXwJQPvogN
GtXKYbZHquzDIediOgT9CKr7EdpxBRR1e1K/mbdvHbDydKQSC2nr7wag6EmMGqRd
Fyx7lqPB3usc0f2NoRlKwOZO/8O1PBbX9PnmJnwqDdiSCqTEz4fr2zAD5L2foByV
iW9TeJJxfmAW3HBdfiqIhaqMoPvI2XXYzEk4+4BoUI4zgXa/BwfrwOCeGFmM+mQZ
uz8dsaeCBV3WRfUUaB4WO5JazXFZgSWaDmKym6RcQTZrJRQPoaOxdbSoszbT5EEa
7FvoeGrHSKqjEgkcN3abn1DoIHvUlEokpXlHaSgbL23QVLZupqVH7ogp3O70CePv
3mAFPennNYt0D9km8eJGGicr1EQvKwu0QpOrRqpmSHORUxn9DltCEYQdA52WfgU5
P5+55fek+tTdbCj82/W9HkKLISyYGxdNaYURgKlBUUb80j6SEX0lvuQOqU+aoRHt
AVHGALp4mQBnEOWGYPSeqWQ7vyi1inmoHYWQcKacJnn/G/eZvtraPoAJhC56F/pc
6Nt1cNAOGFEehLWrjwj+W2iN7f3JY/5Q4GxpBLak29p2wZCUgBwP0UX44P2ImhHt
L2UjsYUJsWT4MZKwdluPhlGHJQOKpTEV7+5RY13H+nRkuSObT5JKRskXz55+fiUO
3rwBIqrYN1vqzEfrkEcHpsFZHCx7/FYp9KzSFbxgO5ErGeExvjrPP1QaubL2UNr/
v764qhXvztmO+Idnhf2/y6/E1FDZQJrscZTRPkM6u29d+5+94ePtleBuigOjdKY0
O/0GzWF6bxRTZQcEuq0tMuVNhR3QP7hgTx9iCh4XtP/sY74wqcSNZgfWGvs2zGby
eMKwmqOftH7mmO7HPTZsWVWt//qNi2QaurY6gc9Q/AfcA35aek3P7HPD+Oa5rJgK
UwHq/ho9q/J3C4IO+xeLwpKCRv9nhuW/8VwVn7TuMV/9mDY8f6V2LZpV/wwW5nHZ
USTLyJPV0nBmeeJaTuyzS8EG3QPlpWS1haTun267oj53WJI1M95g7AJYikp18GKc
WZeg9ywfkg+xPf1G/H/QLHEDJK1cuQrnwNHwhB+Un3jQs8Yj0sHgxNVw09iLwd0M
H32aYVPfGQ9nNItJ9I8P85BmMbjZnkx5ioSRlxwKuGmMHw6I0t/P7DL4Mlr2p5h0
o3vGwauK5MYTYZGWFKZSaqqd89BRTsnV0VZSUmimXp2fXwDcau+Pq+fKa7nfcyZG
Pv2bwp/EOJuyRouVo+lsnjKMf+afRVW2W52yDwnxglOd4HpIMOhN19tLoQw5oiQd
RLDOOXm7sUkAfln8ZjFzWaKIJILFN87ZTzBRPBqf1qvD6qx1U8cgPAH+xYHfX3kd
yFd4ftbtPiP8nWm8JRrQyfCZMCe77fZ5t+9ImqfSczQ3zvxXw/GjKL95IGlllpvZ
Atkx70CuBsl1ni2/PK+IOWRMV8THVsDQTJt3+zAV4AawPSc+phD27tsM/q/mV1kM
RGCBDNekh3cCamLdkKc+Tu0sOPwz7fiK2AL2najkLmnp6lOPacDll9d3OVo3BtCx
LE/M+oIzMv1jDlxBHfqWKcgCNxrnNieoM0xmyaShZVbrlp0pQtYDqsx5cMzKsfY7
P/Pa1ZPJz35c35QHMpmPhXbQAWWL+iPzWUk8ALKp9tqw86Nc2KNtLvkRxePozhj8
OltXMbs+lKLWLNgaFisoVjjB0uEaGiyVU87lXRa2NUXyFjBQPk+r/l+41fQ7N8hq
JgbT2cuU6vW5DY1rL/HQJkRDutji1v6HhdyXDlm8w00W24p/I7EcAz5xwjoUxt8L
mbJpIkTCvfXIiQh9lmIALXEaaIua5/T3Cy0lelJu1YP6mqzFE29gcC8CQ5RxPTXt
tIyq9/Efv7AynWTspMf6OjSWEYSUZBxe+v1c3pc9k015lYiluVsQlgQZAc2b4dVQ
v0KVlGPmOOZWlznXxguLgNVSMfJtJzwoKgvTcZIvrykNMfLLhRP+wWezlzVbCxAQ
gZ6QuQYA/Vi8TNTqj15Ezlk7PyFYSllHD1Xv7V06P1Mi73cHqZ3OiTiunuDHv6XK
4D+24T9Kox9zScac+C09Sg==
`pragma protect end_protected
