// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:52 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
bB6iTk4yqg0lhMxXSjZjT4s3Ju/DHaXX3i7foqPxvvHaH/0h3qZTAxYzf24tJ82G
qF+s6IGY5qkM0zkCvk/b/Hyw2p2FvGouuqE97yokRstp6iXoxya10MX26o9MAn/e
bQwLB8NUtSMmKKfF720/B+rsq597E09LpckSn21UxDc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5376)
mPEr3PySL9z4rW+eBsg7OnjQ3FWZW+vYs2EwX2XjXzYefn+ZzAPZOqmIW0odenkI
xRS2tHIiJ5T/DQ8MHOE/IrtmmW/JLstXusL81wtoAEI47G/2Ro7FnYSUB7tqvfGv
+FcqS+i+T7EMfW/AONDNJDWxDVUKZn0Ma9kpVshbB1qEu1FlAgVj7d6KA2QnmRmv
eAiPj8BH2RdIzMyUwQ2XpI6rw9b6pG87elb5kOSJs0gs6KHHRhNGHlR9rH4VuG9l
C0isQXSy7XgZltcbBK/ALWzm/Did51ZwfL7kvptZ/8WmsmyuURZh/CGWklo/oUDY
vbCErIrgxT2/fvKFnudg0YYFook3LG1agj/5SrbbNpjJbwc5QZhXuu8RxItdG+jS
s9O3VmSoZvNi1WOo1aP/WqiZ1QCjCrOL6JxfLGRF3DMmK3QqRIe+odaB1Se63Fk8
f/RmreIUwAiQ1BZ0/XHKHAx/tLrMs6Th7OUl5Zuy+3328uEMznnH15tT1O4GOjcm
2CL9vDFMOCSogwSGVufQdTiv8yvwD+MhXBgZ9almVTNb61CJIZDouMk6iiWhJJgB
5syR7LXjzcTE5BaFnSMChIrfBfSFb4lWYTZL3eneyqRWFBQXeUlVqtoCKwuexQLZ
8xYF+KztmMOmZiLIYa6J71tsL6t+foiJHux3ML7F+GDWmqDdo4JjFDSkTrAQ9OZZ
QI9JeIlxELINDfh1OfQJLj9PS30NKbP0upTiRI1VAsrPTqOeudkenD7jHodpyriV
rhs2frEiVRw6nG6r3ZQYVEwNJtIW43bcexYOwdVYdoMjB0bpXOOFiakYfE7lbQCl
AHHVLb+aEd+87EERzrChg/zzNqQbFkoSvwKpU94DSsv002N13R5BRu16joJmhQb+
RaIqzQNibupIup7Z66ywx02Lsv9ibXqk81viMgwDoflU7RAGAfAprtb7zYNGilLE
r52J010PZj3GtZ4y2NbKV/JPfXviwIVfOyFY5rXYXiHalbm9dI70krlNqCTB1C2d
2tkkYe9GZy2WnDcYgCjvyTgBPmiK5w1NgFJ2HE/N0aXHKzylabN945gfB3fSd1b2
EOiXd/S0s++z6oOAJA4MUi7z5ECPxC3HDDjOyYjujRHmv4BxItqAdOX/9l44bCAs
nCxHoNSube+Cpb4gCLG+OdsjaPI1GSv3QiaQp9Exz/YXImOySJKQGKs1ijgN03hZ
yBMo7q11UkHdeTUnYaeikKdf5gWdR5udEWPF1mXqfPtuRgylHCcENyyc3QczKOFm
XQ4RPdSmmw6eiaqrmgf0rBaeFmF/DqxlTOcFtNNKBPfOsedxSo8h0KOHVK8iG4Hc
U/ZFrLw/AKH8xnzTOX7pK9vqXgt5RT6LtJRP6hJJjUiTIIsSZhsGvDMaP3DMjYeE
EO3js8f3NEXnUSr3BFMxVy0ZMz5vVVN3XegjC0gccIUS8v4T8n6Fp0YZRiTVgOu2
dNX3Hmsv5FNBwP+ZcB61Oefv0yOpdC6VG9YmbmFlNEr2KRCa7TMPNXscFvcjhPSw
eBHvty3lb7Bsgz2LukT4/5mhmAKmqevvjeTBhY40QtHseDfNwL9MQ7F6X0pj/WJp
IA7Ukrs0b5yukDg2nArxap54JZmroN9HYd9iPLYFtIzld7XNnsyUsPAhXIW5vEjU
P41WXIT52CSK5YXZQMR9O2uudi8GfqsdGrS7coR9WeJ0uxp8pFFrfo7Qp6Z0t8+G
NPB4peVhJe8SPhDBpxiUnzOiOyC9aC/dADYVHp0w3TrtAPj9XvQSY8To7IY817D9
/ymB1LwK8K4GAy1Uy4E/Ck5HLlMnMSnTF3FMctoiKVXtZxox8/q3xsOe8U8vzf/M
qjlLts895G2xt2J+F6EmjnhQ6peKK+iu6ASvQlPseCln0xCHU28TZZwdNxEn3Pqx
dRX78HXvwbLQinI/dExHoC64yMcPK82fadwQhX+3VAQW+hwpq4CBc74rokyZZaTx
I/4DA1229Pyj2/xApi1G6q3FrEuk89MUrQqEtfnkOTuVJvqYkeBEJjMifDG73/oG
E7ijnns1ex0J4quE+fihtll0Rlk8KY68osc5ZqRJUCCaNTjxJeQu3OHLPW2t8VYD
XtdfO4S+6dvTvkbSYSb1OBDFpc2NcJILG3gtPfruVPtdn7IGkruh9Flpfhf1zRIn
zQRDQk9y21xabpNRUctPYPD5OOEd0+dz27Upa917TXq6L2h9+g/Ap2y5HyRMmkDx
6E4+KzQJ3WtaOfKBTt8ofVjRKwZ/fNrcxI7cqr8RqLKOZdKsL9Ni14sVOgsIEtJt
Vvy9Z0VCo8rkfdFUAYuXQxKjabiygXidCZen+X4NtrkcdNx3pTBlmOI7aiDJfjnK
/mJUSHTv2Jf754rsRYuQ6JUPVdL7CSIls9QjbE2qMhn3GZ2VXJMFPg9iedyKk5gd
h4chNYm7acVGBpvXiVSQxcQdU6yuWdBpoC2zEkdGThY2xTihleWPzx+2Fba1g5zz
8agZrVuQnm8v8trIsoy2OyckqD3cqQRcUmfWkcN7f6gy+TM8Eu3cIm/pKwiDWY+g
uijl38iMF+9h/hYxVAmGFNoIO340sVGLF2SyYdO4N+oxwaL5rrzs7jXjaRMncw8G
qzYSVhPjTNqYfVASfdz9MBkF3OzJMx5XwjQaedHHIvEvnMtrayepyeZG3dE5x8Ad
gq1wYuVNgnyUHHPbS4HF13RA2QmCflrAPB4rnF7hW6mMcvAvmQOQx2mPHEThcdGF
C3hoSB0DGZYtJg/QVgNLZYKhmS+WvwJrJ8Jh4K5uXj8uupsWt9hh2ygU0NrFhzSA
kGNrfuSta6JPUcaoc1+2SBMiPTZC8qaAn/wjLMuISQ4g4M/R/Kuo1u9SWZqU6Yb3
tLQ1VKs/PehTG2mMHDh2BT/N2aRUa3BwITsY0t7PmOU2yK+GxKNGXEdt0bjIY2xP
nEpk1Ki5v/XfNH9hVeYUVxJMQkPaNgKiGMeAM1FB12kCPD2QNAvrhTI/gz6T0NMQ
+31XCYxo0cNbRSdgVpjfc17AIXkXaG/p8IV1I+9PS1a2JblXeUFb49WWJ1cAFXOT
2Ckjt1PshoXAPWSAhdQEdIb3aivZR2PA9SMHY9Y34FRnyL/LwKGD38UExq4H1TI0
3/Ui0QhZbS+bhZuMdiolRXQDbGTfLrI31QR+7PQwuxJO9A7+164HeAdeprvpXT14
rSXAT1y4iYwS1Y3tC8VHMLFG1O7fMiUBb2fH7DZNs4d/8I+lGUUGWkYitZnBFA4a
MrtnGdrhLCHsGWEMNy1zy+fwkwIWviugAbk3x3IG8ZoLm21lVwFDVhfguXQgPgom
2eDa9mGaBmQSGOWVSfwRbMfeYy9vN86VmiCldAMv41IjSVDirCML16rx9uTlSYKE
mn/umXwIafT3rhMyR/XGccrPlBBnIDRLz+cj/PKT04LEFl30TPWvE9atCPIuYm+R
RZWDyVVWbzvJeO3eTnXPUyppnsMpGD+3yTYFIXWMRD1pqtmTRI/NbLjPdorXFrXi
vJJmG2/P3LijeEbPZmaeRpZKoTKtykztXMPatY9JqVgyoLU0H6gJLVlfTZoWu4TL
Uw0i7/Fkg6OTNNvT+khZvRpOzF4g4xNqwjNTCiDortzO3Ntv1Eoa6v4R2IVJlGrq
cZZ44GJPw8K/fH47VZPJ0hEQ70Oykn7W2unA/tUbAdtBW/rLoriGzI/MJpm3gsZV
F4Hx0oTHU5oHl41uWImpKGctPtO+vZUMC0Gt0sfbcZFEJ4JnYmzDdlX+A2WF16zY
DL7OadXuseRhL3xP8saguJtcYcmvOSHVbGeCFXTLC4VIx3B3hlsZfbhWZpWW45IN
1ohtJxCDL+eMvUWSuC8//wrWd9ilDnABwPbwtRZuFKqwmjrZd6R4rD0TGBg/HwGp
sOWitG3a81ehjmbQ+2q4I+DHMw5TkuJx3tcGS/7l/XWAiJkfWtxFvHuZO38UBAxU
3/mPUuKzgwm1zOcO/7NkEBwofjnHdUbj1+Jms9s3JZH/LP1/Y0eY8q0ybJ6K9Hta
CeYrAbySKy6j/q2NGxwXmQnkUXWyp91oeAlLksVYulZk55QaO3biyAcMucInbKXl
+OVSVRfuL0lciG3B0B6v9z/xIk7eIDg4j5wfxFAS0j52BLpub9JE2qkk/nl7TXOD
nRuGXoEOHEb+WYRonOdT+sZ0YkVuyaXFTKF9nXy6wK0PzrP/apQqAYnbcb2kKcG9
4qvnieCj0PU8Z1Cax+sAVwFa5vd3ZkFU59ITknU+hRXze/ggD/3/Dl+9U/yd89Ov
jp1an32DwTQz2v4PHwDrQ96NHJRGWFaSzySg1AnVC0WzZfPI2xnfqntiMMl6VGBy
rCqP+4hvxh4VJujfP+ys8CA1hA6voGMm+72MQfiM0iBWZ+8Yb00ixv74Iv6tt5hG
MzizsT7rSnsf1WSiE8Zcv0D/JSlIv6rOfm4uvxZoGSwcUfA7vM+aBes5XX75lK6L
VDGE/k6JtR993Ts1m5oYDTtdQU0W0qkqRTS5PKd5VenIyPTbjEw9QJuM3ZoYGznT
AkoRVrentq7dMcYOhN1+0+r4W07vqPQ2kzqz7NsYRWFRWFJ5wU2jBYWAdAHyf1wK
yABgJicZNbpko8Ph7qhkBA7IC2X2yzvds4ZGj1Djuetbj4OTjKwqy1/Gz1mnLHmI
2shuy7qb/pCAuranmA5YmyNVlzpaE5vTQHinuZP0JpNer5Uz5BAB800NNhAkjFUN
oLlp4Jdpsb3U+JYawX0g0bkhNoe1u7NSKqwBsttnNvGAayltj+lFbT2M8qwGr3Gh
79CFFwCnXLtSNMZ6fmpqnjAhWtTDXrrdkIb0ypWBoGHM82JT8sCiXRMdE+CyLzxb
O978uOFaNbJz+VvWJxDsTmuFUjDLmPRjF4w32aJYeiHQdGSG1N7EFiwq81RY8I1W
46YmkcPPK8rTDQh/yg6euu3c94hrfZZYhCbLZLJrEJc4hsGd8kC3rDbZmn+QF1iI
B5omLSDfW3xAQVLPlVOLDZlmuJOjpIxdXOcISEzLKA5ijKHjpwuxd+LqnBxNf6ee
LosTHNeYISGFzeppwwYE7X46VuE/0lbuantvhCl8Y667BGL44PZmURgpMs5LUM9A
/8sWwKMObqwTNcWrKrpeZZnP0hR8WT9f2SJH9cuJytZQG0bnYCb6lLqhInYuQnBh
43oB4G9m3UiRr8V+0vxFSVEf4PJMKz63rJRiSURCLY+vzjOjcmMBcPVSt4En1oG9
idFN9ExLBxlwbKx+Mkf99QMGerdnhcT0KrXZNBiJU9eat+AIIrWuGwHuJnkfYbkM
Palb1i07ReAQbjiV/osrfFm1H3DxCHQZCDNCempZCo6a7ZRtaGIlQoF6pqbWZ5br
GVZGNLHtYF5BskqWa5T7e7dPu/Oe8vMEjMnQNZU4dAYDvELeI/Lif9h3qNcPeSkd
0jLY7waUyYiGiZmzZNTPVQnMHEPDOs3g4QbhJsxQu5Y486I9iR8ZKlA9ztzOJlkr
MqNTUBB5CIUSivE0kmkInCqtuBn+1H4tXnImN6SBJJifK1nNCB/YwnrZrpBVfykA
JqgHP1BIOxCFQ7AQZwbk4Em0MSCb7KL+LyqYUERayuHo+NmR02IiihOAqBuGraNV
s42PXA+vdOzY9aTgXUlsJhpPFQ7oRdPNHSGmioq1so/8SYyhVucWfvbuQ9vPopsP
WW5mWlkQjAQM+7VKjJDyYOI5kyOLhzvW0uIYHqxpYbNIlbYiD5ArhbGf8Y8Xum3Y
L0hRP5LEApLKxF7rgmiHre+f48hYKEtcOBUIq4vSfmdBO8U8orjEMfmVljzOHTzA
HxblCO/fxtVDZJzT/mevq47hEwLuteJ0mPyoV0NNWdLJ3gdHHTnodlAHNdvp6JKU
nRMbFwKIIw2umJ916tbR5+2bmf+ESw7b813q36ZyoG0MZdo+aUA7j6NPg6LnOXAE
QnkyoRQAGXpKIY05VY4hdRvOIVmMJnoPcS5HQyiAgUqm4VbEXZWXJ2ioQP06R3GN
Wkpk2cKLD2w2bFmaAzF+QvpIHcBicR52j4hRjAY6djqAzIMKoCtIIh++rusOygmS
rwNhAisQvxNFDnYe1SvZTKOnF8lg0B5vYsnbqJnd4ulNuJAtGOzqvk9lI/drwoHn
PMguIDFxvFDmVai3yIdTKa1iOAakSIEuHStOQ53mFHILESUHL8Aebq3VNoO9z+jJ
pjNyWWz1gZTl5Bj0Pmd+YllrAuQA8WfMuexP/Qr4fLHtJJKGnmBw2myYoTy+T2E3
kXrZgUFTlAShIBpJltnQLFpTuRD6pN0yD9fCwlDjeGo9gDUHambsEkKNrgmBh2Nr
K3WzgSUe8KQ1HN/8dnvwV2e9lgSL5e88MJzfePRugVLkrwv45OE0r1EBFDsnZih3
OAcbjWW0rckl3GBOTFi9jWkgG+5tPuARXnZeCTcGGg92MTFTdX6jn/bjo8LhnIiZ
hBVstbzQ58hay4boaETq7GbJvFeAb3IHb/EObJxxdp0UyJnIDnWQ9P49gpGKA9PN
wyEGEDpDRrNYZXmYSsm/xBcwp2fknGWXWKYqM8xCuRHZDNDhj8hRRV2EKwaO4F6b
zxHTqTWaesUP9bfy9PJmVMGwvan9SPtkbbSg4lo8MnK8ZyViYK43EDyMFH8ZmjAc
eiR8L3AQWZyagcqLuEULcCVeQtuUG517xgd0ZbvSxpbK3rYK3V5sGZA9NV5mrd7Y
1O/F2/XW/XIDTN1kTDQJ64FQ+Bm2V8Be3Y3VwsRvXckHybSn6dPNwycOvVYnzDk3
AaAHzcmkKx7Yo7ilgIpZvOnR1TSxvxGE+7ryCUGKzpy1mkFaChNgThhvH1ezInnd
kyzOd7Xwr0b6jchI4YFVmZBHcs9HOFQzrws8GE4VSR9fTYn+yImTl7pHBIQZiQ0X
G76bjyAnmYxLGwLs9pjpbsHC/Hu1y747dZDWUCnozBJ77WtOXwO0sKoqsDb2j22q
rjh7d3OGMBtVBmxpmZX/jq+u6Et1nAcLH4IhRjcgMPojDesI1Fy9ySjvufpcKMoj
J5TtoFX5cVwuFtfhYW9VpBULKcV9s0fbAT0Yl5Aql0V7yiQTgmKdRD8qlMiGrYSd
tS1bgpnyOhvpxxRjhKs1ygvt+LvMK1KdMWc3ueuodughmH7Y4lQDisIZ0honXdHO
`pragma protect end_protected
