// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
6XHaOPLEBhQbsltTyierGkwjwnSA10PhQBaW80ARhjiCyfXInSPOhiJKs7PegyQE
Tz+GTVsjQaLP5VsR1DX3xrCbruzflc5NfzrsitNJLs9p48oTcNDcro+rN6vjP5lk
d44kvhbnQapkW2LGaQjcPuC+q8DtOa88L5JOYCFg7h4zLXxJHw+QyQ==
//pragma protect end_key_block
//pragma protect digest_block
aJn8/zy/ZzyY4LuWWgWffOYnocg=
//pragma protect end_digest_block
//pragma protect data_block
bZo3OBr+TLM7TJJfIfcefBjLzdGty+yWBs35gcQ+K4f/oyA5zZMy4Fqaqk6l+fR5
Ky7WbrxiD/eN/035DwUhTRfpE4pFaGc/f4wXKdBlEDpit9pW/giqtRzoVfGwvIIv
DYHJPmVeHT7sPOgw2siliD4efCWuK3oGi4O0/tj7LmfbgSmgy0GTUzxq5TlprKMf
GIUlOKSba/kEzaxTz/JPdHK9NXxNLCWScw58czL0j5B99kpKdQUySDwpps3txs7X
CRsTSli9dl1wWpm1Dex/ljknUzCkZxqqwI5/YLbDVlM7yXZjCeNzICmnFcP+39H7
/YkiyLG4KDl4K7NhIELT6w22UK0LX4HoPBQ/dgCWQwPLlkAPYWugOSCurEC+556x
wuEQN3T0qcTdK9d/1YwczskxjvrJdX9QkyJqhwfYl0ixYzQWG1UPa+Lkqs05FLq2
hXk7eZk35h1OEd70zL/DYiSncjI++bZ1LbdPp02bsz0U0SREBBjY9LmSucDz7b99
gFRkjfvwZuqBGtVic9wDJ6qQG5a8MptgkI0RQgqxNQLIofJNfRunK2x41ETyIhP8
goujIJFY1maIpvAapvzqw+CF22nUjZsNZrXbug+PW47bxFzbOAtdpsKK9swyphpt
noOugzBXoWU0ziBaUx6rDltDETFp3Dn7Jgc2M9KkW3cGXE5mn1/PomxBNdPAeaQu
65c3zQg94JvFLb34wl7Hq43Jqw26D62MtaJuiYi8sNUsfy4W+q/Pe7uytXpqaAgj
b2prS6YFnsJVDrbtEziCxAMnOrHzzzTnNG+pxZ8yCq60kAZ6Ih08UlNuGxsFzAbZ
guJkgfYFgOtzD/XhrPNPYwGKCgeJGo18wL1yzIfQFCbHK9SS8fE6NQUKUw9CNDuj
Fe2sBd+sbhaOm055AtE/VhEa5UNbyHEtUJtdtzFxSkAu25Ywn1Q+IK8OTXAQdwEM
eKq0mE4uIfro5UOdfQmlOrIHim/vIq3CtjYmtT59P38qoW9Z0Vd9OSSpt56b/4mP
7ixr973r5kdiJwsWqroXpU55f1OkfLn0CBkoSAjkJ3ekZe+/rCiD1arp7iwS/lKR
FBsi8kSfm+WnkqQ3KYUiWad4Gy3puOLlaYO+ZSPTkhd8N3wdi44Ta1864oaNctfO
diDP7JYxyC3AIJ3I0l7LF1N81teRlW4tFvPlHP5EG7QLZMpQi3blw5mj6F1aeOdT
PFHwabJidyLsDtRsunBuOnmpp3X9GxDTKwQDUmG8hVhYLaZWiz90xsBVI1WoR3ag
usXQrKQ6u+WTMV/Dkbk/Qv5Az3tKmA9In8rxAB0MPHVTPRp38vuV07qB+yFm6/+/
TDqcM5NJa6l68riU+k8WPffAT1exSR/4j3RxGxAZwAOT1OmN74ljB/Mxl2Ko4JyJ
RbzHxheKGFermqduo4ddBYdj1PIJiXnTFPife35OmwwXwqlm+1EOfsAJh88uhvkE
2kW4NdnNormC3xr+4hpyrUKcBNXiI86Ypq8cdybE7teMOlHD+5HQ+G73q9d9r2kR
7qn4ZUZaZPGIWA/tdtwLfrwADcHl6/Fxm95SAGciXGJwgevTK5Y4wptIdhM/Fc3w
wFBgUUSStmHFDiJD0G/DqHtOpdOUvH3yGOT8M3etrTlzSCROkABjRbyGb+WlXF+Y
5By/+T8UGuCcJBlK6xUlOueeyv4VFnyhxbdY7m+wB0Drk09SHJfA91hvBqaGAnyC
vfKoLrkULifg7Ei1RaxMqNZcUpjZSuAp9/5Hu0rycMARn13+ChOPT1HB2VNmE3y7
u1jKpWM4NRuzxMsub4LVEKPh56OJbEyeua2UtJM0lnBJoz2NsMtqWcvbo5/qYvFQ
MACAwc3c8c49QD0/HWQ4xboGdWiP4LnlVRoagSFlA3ydbaI+cDgQl8w3+Xi/T98/
DM5uBmQaw++PArbIEe6raLucOLEXQcGnvKDxM7wD5Mmp7dFU8yiV7f5spicWcgSA
YP1ePmUtcu7ZYazPxqAxMrsIm6W0gpcyA+NmMkLc2KfMxxoaUseHTiUIBqXQz1I8
RlSNIypmJO9t03otmJCX6IlSlEBBnn89Rbqbpr1MejM2KPI2+hFSyvjHZCwuTNdD
cvJS3Zw17b/UWppkx3mHMEJpE0ODE6YcADP2C0Ss4DUU+6IufOo6UyyUsSzYFVwe
Fa12YTVVTcxY/j5e4dilm+/Xvc7FWrfr5pOzJFxkggPh3qXIvv2DBLI7+sm8oE3m
hXDdpmavCpSNQGhTiAn2EbIcG3ALU2AoN626GdJaYdFyTNSzrL85yfXdXwgR2L61
P542D8zAH9fnLJJuZvxR41iMunpaveF7G8jx1cpYCfLxRbo5kugFLniJZxTtpmfp
yEoekM2ZgnSP1dG/BHMIiqkMNzZrc7oxczsbzUbIjCL5aEDgYbJ04KTCvWoyNoxY
U5EOZpOqrimiRxx2OpBfZx9IQqzGmx0sEMcK3FEKlBNYoh4KsHbG7NWtdgQAW2Js
RyTbq1pkNbzfUTxMFTl5mRFXvAAjuPWmI2XFI2W3ASKvhpDBFWYaQTicj9i6HJm7
YI4gs4sh7YiEmNI7mypsnQD208L5SHoT0Q2+ySfmUR61/BjlBRTjg95qOHXirtOG
YQcspmEZdNwK2z7l2BDy4fj/ot/UQoB8kVHeugnLB2VDKNU8gmy9H4Jd1XrZNY7M
c2ON350peJOUanjnUpSD8yTCdpAtaCPPJUrVs/03m0tZkDBYfEYgcw6LCIdeDRhL
SUGfsdjeOePJHQXHTkn5NpjKiCkCJIsoQ9NPqDr8v6TVGRxl0jTprr40uNshJVT3
HMDlZy5Q1k6CrRfz9NqT2gbM06hy6b0D3K7Q33ZUj3EM0f674fDTx5ztjWHEdsQ5
x29+WiCu+fn8C/y3arpbiwM9UQvatQl0dZWYaGip/0s0xNkjLUEj0c+FT4LgVdYl
z1W+532h656Yik5qLp/6gHyJi0aecOL51Kh6uED3cuoiivQnqEdIcbLD3quCGO3Q
2ShD6aC/kUaMyrJkBkWYuFygunYlcVS4z5Kv0aKLRY/cHR8Tfd2ZfpcmjgXnIDQn
GUqM7qoXosfucdASO0qxDsUALdvzaRa1G7dg5qBFJjU4wo/XtrULKNtpUNaR0be7
JtVy9dLFM92Ugcxnh4La/+pP6TQOtjBOu/sFXNejl9rppIBA07Tu5U+Cn2IuhQ8f
8R97lOhzvre8iip2bpvx66/0xlVZ2BOi9yskqPM7zEE5tyfyun8SnNVP+IUbW73N
mNLnurQ1GcANS6g9QBXc1mzpAeMsd9vRKtayIsSnl8YC1UU5bizJS7YoIYrM2RKz
zPSpiJzAEAmXMQ3aUiQfJHgZuIzhcq5LbEnPI9f/gZbfU/1mG/r8UO5qklI6GMGJ
eD9O4Y9la2QjG+tXHV4ghxYfzm5z11RKqNJQlcvBpJrYPy4n/tvDKzcdtCai8w7o
lmB8Jp5/kC0dWgTyRiRCnBEKsnuGc8Mq2f63OXVZr29GghWOq+K4HZUT6TUIGTT5
3gR6Lttk/5ubcRqsVxvCQPOqufDVqrAN+yMjjDmQJO5bMvYU3r1HjbwiakWSAszo
jHGTJsD7kULODsSNSTUyXwbysJS6QoJ3LZXzhxsz0Nfbj+OrrsV3YgKV5fmCuH7r
cqp8DrExuiRwvrMi8B+XuQnspCebketCsJWlRnG48fjjWUUVbSNTctGC0V3vowfK
oBEdQYVlUrhRepmJmfyaC/U+4XnpUgXBYc5ivvHu4KZLzCsgeKPjgusCRj5DPwMp
m4AQI67jifMJt6NeZt/HK7+Ryx5jU1OGhEDlNXrGw5UA0jJeCS1rnOMaXWlVDtjG
tcdcarh9OaH8gnO471G4txEb6IEj8aZWbIGlNVeWd05DIEf6hZXBhYXNHs2hH2jk
xBRrtCTtBrWH+8aMW46wQYSNuJg1sQ8WQqt9QNxt0U1ziYtXqslNkxIBgvZBlIq8
kVRTKuN3TdycAlDjq3U8WOu4CdveNE0dNC/o2fW+/GIl6URmWBMNIXKJqN3G1WhC
7Or1d1wY7k6cBRhh2Ox9J3xonvmeN1zSqTDwvwIxe2OVbFhJmtXMEp+H4LBPNuup
mdIkZwEdmcYhGIySxR/RgnPIy8ksMtNDyFbVT3Ige0SMV6ML5X12b2qoq742npgw
K6+a6h18lf+b5qVZnXfrU36WtFKuWhIXnxI/FWNzadvmzR3EYKviF3iNvCubI+3R
Z7Wt2EBvRwy2vOw4DQRkeuEpejM1UPB+UBhIj0N/ENcLUv00ECdp2gqJH/Yp+lpk
5pa6j1SWbcHsoKnYmluriZUyDvuy8424C3/ko+uMBDLiLZmy9dD+pk/kdoMOfsN0
BJAU+RI0AZ2lgNjun71JPArNFwPyhuTJrjs0O/lw4f8FjsdvTe84e8TlU4iEEpHZ
NAbx/ZmOi2IC3fR8HfCQMJ4EylyY3/ioKJy3zTc8J2L/+J62gfGzwSnfqIm5M8X3
vcI2Kzkte6gT0ZMAxL+8rrm2tvMkrstBD6c3hwOUmeTgaTLROBxQ1VlaF35h4pg3
86bIuxYTCKDHwUZhT2Pk5Os/N2uP5l2V6gxmUSqe8y5TKZljiKHEh5QKCLzfa0M1
feyNDui1qUkP8L2dObN6Ba4FZsGe7Md373ggHSd39wua8/0fpuq6c37GJHQQw+yr
IDGUj9j96Cn1HgeluJ1B+Xnvck18uWGFKhhkhebgdkg77HmS9HVeW4KQb+LDRfjj
+H95oGiazHbnzcwkSw7xpUEYr3y9gXGwr/mZOFCX7jvCFWQXGbfJihxmPuMmIqWU
0W3bUMChQf5aoLhTjr6tTK23116FdOA5IWiDUWSgz+mONjDluDcoI7rhKzG5HHfL
wQncCgA3+f7QvXcResI4Rjt+RgGoaOhn6wT7e/BfGJsHEt+YVHJ79W2MGW9Eh8hs
GkqF3svhFzzvzgHVf7zwh/OChlk7t7miXkVx5PSuJPl1UuO53fziWBNjs/fgO4sz
t5Gcpz3mZN+DwWLlSmasjxfRLYulXPluNRfIzfNfLOI54qeaxuKs4Yfn25YMl7rZ
zRJ+SnrB6GI7w+EWPJp5ew3Pmyk00+MVa206Q9BE00UA6f//iCQJetnv0ZwAB1Nx
TKVKwaEBm48uzjTs/sxlm0sUog5ROVomC7jf+WnlwMt2Ny4i9xurIy2f/+IyuOe4
2i9E7jSiQfKp+f03kS6PdV7vI7/6+iJLnZjviE5g1RlMfbRaDHmnDviOz2VLnPsy
xVFqrdLp6LwD1KEI+tjj9Yh3RzOz9TQOn4cWTWi+qp9j+0WjmdUpuqbA85Qy5Dxc
GNlC6NxNyZlzeBe2RN6U4OG6jdL7vDB+RfB7EqqU2S1AosKAdVK6J3ioN4YvvJhJ
S3wt/WF3FErZotix7KIHeunhBQ30gkynfrbsoKE6Y79xWBypdflE1jS1k0X3yWp4
L6wDsth8O5+JOmR7vhrjMWdNs2Ptx2+QYiYAlcERqIWHhCSt0uzKe82lbRx/JTgB
xhH6m8IxgKQizy0e3G/5/NeBXmtyfp4RKIY4YVlbeWOAPQ2AK4f9hnqODWdMQnZ9
w30PgEbs+3xzsouK61IpesPnNJg4+zU3x/a481goVqoSiyzId5Ap2hRD8yilQ+Tp
LDbj10iO0uvcZztMJlVmnfQxblMU6Z270Yjjk1Vaghxa/FZj7MOftt5NMEcaIVGf
OPSFtV0XsXmiIShk4OdoUY9Os5Uhz9uOezzYi6T21MCsHa163J4M6TvDfratfrsI
LaWm46X7nxh4WC50P6/qwAhvRcvgIS/lh8G1Au/U9qzsi0qRsLsx6letum8hq3id
EP+SzIWn9BCv0zL0SD1om0HnJMkEOewQxKwF2De+uGLwIGP1PhB1yG6dFWFHQBmU
5jXXhyhYsYIoYRTBlzenEeH4XQ2649XFRCSYURsIcM0nvbt3ty1CzSGs53cWStnH
tOa8eM1HMOscCHv4yecfhea2ic9zcIXIb8x5k4z4xsa1I9sqywBaIth0l7MZKXYi
7p4uh7oidLW5zgSy+4rYMqNOooNuC99GEWau4OJ9DkkQdOH+W5z4VmTPOEzNOFUM
RuNlFiwOYvzYjSN+XofexuzT8IBfqcjia9qWRxUZxoXT/pKIiTpGA04zbErrP4za
AeaWGP4EqLcUqkbVeMz3Mb+1hRITdtVUMCq6rgf1aDA8ppXBmx88g6BIELyk4KQC
Rd6nri2Ayj7iQnoYR1AV5QO8xKDMFHpEncqKpzV9bWPr+3FmVqOYFve6aVLoz95j
Rbq+t9PXrxVonUuwZBmmZ92nKGdFDg54tZRmPpR1afP3Q+OWrmju8hoDrsByH96n
Mz34BZn/X8x5ZznJ5GKr4kT80SslydCv7f2u+0g0fzYdgwhkk7r19zJY5lDgN7oG
t/9neecMAE7Ru+XFaDlJfLwdj/IADcSpBftTlAsJxSLzaoa1F/MfK4oUpyBqdZi3
U3zx/gXn9RG52ZPfTRn9Yfvi7813/XBTltPcCr0Nj+E36JRNh9dNEQLeVyDbMh1j
C9P8p3vk8HSLLqogqjys7p67Mq9wugeu1SSEjl6ccw1rAeNdGUQvQTXLuuHnElJW
p9H5DDnoPc/w3BgJaHDu7Y38IpW/QPfWerQYNqCq5wAvaPm5LRv3j7z/Ir7bkoxN
mfE+LVt2VwamCqlCydkRN0pZc2FXt8zM6Wt9AdLQZrOs7mmV1qsrH2g1nUkbPOjB
W7IZuUlD0egmOtYwlluGVsVyKNU2JQxlQdILyL89CCybD5u9ckndyuAKAW4dNpLo
8mS/aTYpV85Wlr2D/0Jcw3M97DZ/czph7Oz7A+R9/JtEzaNEp8+3yVoFrJ4tNZ6+
+VwOkO8U7eaKGI+qJApabsHqgmJqwJ9DWgcMSLjO4stuik/gACFJkOuSNKQFwpCk
nxPs9Bm2OxTHKKWtmxgHXZcp13F044TEhvr2ekId7AVAdm5h7IdFXkUn39d/Kxh/
8XNUBg0hZUHXnCvYACOkSGcat4SgMHwBtFCbBteHeqI0CsjNqyYvUN6WYb8LPib6
DmGB/np49Ta1x5VI8oigQnoFwWuL9vU350W+ocUNIoPshB7V+usKE7Wz395W9M+S
NhsRa8G2AP4ZKiwzXvMvlE1O2fKX/m+sRV6iVwCPbDCfKsBl37OLWntPUd3rAmLT
i8vO1WTA3WDMhf/ROk1HbvqSky1BRMSKgqM182wzN2m1XcwhRM+DctIhTDvkOCF6
g8ktxze23A/UYfg4fQB3JwpNSbuZnPppTrzmBFBAVpjEjoNNn/o1pw+MuiRY5ZSw
Jy30yLk8CGoawn3jEuJa6Iw+2PtqU6N3XR6o1TxIXqd+ncIOZtsnj26uPjb76XsI
MmUQm2YAmFL+TVhjE/RlCma7bX6jFNtiGSPBmJF78QNDB9meMyUPmcVrEHa9/R0p
tfHqZx6L04QBVq+KVl0Y0TzOT86TJL+Ezt0pAyRyP6Z7D34YZUES8wrVm7YAv6YW
SkcV2c8xNbLTwyGMTCeA+9rAubf9BcQon1c8CWVFb+2DIp+g2s5Vazv1A4JzG/x5
toszd0bj4ZnDf5GeIZu3H8tz4e0VHfFz7B1/7DGfadWE8bRW8J7xRM+YD/Wu598Q
kby9Qd0hS16Sk5XMNYpdXl3fR/L6z1gEeovFm5nrVi+pJO/0X7PqCftyuBAXtNs8
gLUYN6ojW7qqJ/7gmXgkMuyF200e/3pBxOZuPqsfqWBN2iVDK4zPGtIbGjtyvHwH
VQbyHN1FkIJJOWJh3QxwtgWzY6eXEV1QnLYSqWbhgndTZaVCOSdJVj0tXT8oSD86
SoPx/yBAoSKuvFzF+NPs43anxz1y35mxLqJEl3pTx94aiQHxvEJWFM75J316ECij
SqweJAzkLVQnT+N6UwJChPAJ3Wxed3djOggN1LukMPhDpRlz+je8dz/PxYm1e8Fr
KwUb9u23Ahrb3/dIfMPHvxOqZyHmBNmaQIcgcg/wB7j785yvFhYS0Hq1YifbNZxd
TAzRGbnGdAk6dTYyacNolIQBk3XvRNwpnEpXF+CnGyCTPDxLIsOvPh+obNGdZYiF
jnHYT4we9YN9C3RuJpY8e+cxz4Wnfq/o4G/32XVna8oDNTj/TTSSjcjGuWWe9kpI
UlCjDvk04fQx90CwKMui6WKK4BJYUNvMmbsCR7OIQFcdAc4s+tZ7UHgI6D3GOd9e
C3tUHByQPMBj/ZDwa1jSyPCvfxQCyFxbuTCYXZZR4/s5EbNXUQmE2Ef87I5lG9EY
SXOb/kMtIP3Js3SxOia4jekIyQDJrQNbiUWF8LdgZh4TKv3vjAw2lmojIgMu6Q3R
LnxTJSMzKeXAEbd11AKpb0BcpqXDfm66Ge7wjcUhqehSruFk2yXNTS/YGAidTnrg
wi8JP45bXXDykdwvnBddQ1OSrWj+nWFWxpiAhao4pN/K74VuNRsRaVaIhqExCTjL
gsspY9lTgCLMSF+V3zK7JhU4xUd8ixQUmTcfujtz2F4+/SAIKrXnihXRKUHbiLjq
TqHPhDa82xRDLVoRHAllu8pbFFDTm7yhxU0SyCqNGUGLzqs40h9+8rATGMzd7Y6F
kNpl9XrKRHZSnSJpfOm6r2DaaICDTOGnPFGZL2WDeCiSvGPUs9zxynFJFpYYXwCI
gNS3GXpuXLJyOeSI6ijYsKRT1T3GTi4FIwfVQK1heNLPaR48Pi06CtzMzbAPtgGk
FhFmYwIlVjuiClJd1/CW4bWG6WV5vO52+m0lSfGuPk+hFBH3JjZkYqFRDnrSiKyX
UIOAWusRvGTMscund5Ai4J8D91Xprxm7M6ETFjtERmuXbivUfFxHf+KLGw6KRzTi
Jhq4FKF+jH0qMwiAZOFz+bLURlIUmDupmL0raFWlkuTpMFn/Pqs2GI9LTUydSbIr
oqiHlRIQ/7lpvT0OapLpQo8FxlEXg5/bcFb9QFhITIZVMmlaWwY3yf3Pp0Z+OaxY
GQ74ayHkdVm3JFhZM3mJLeFLmXWuLLStzETSdfWvZphfIyeqrJBXKkjtXTTr+ZR0
8HBH44zoiwRXK23mLHAVJbueuQQWy1U211dVc0hQean0qlks4DrHgfVPCaKkE49a
pQHLFufS7+jY3nCoGDWl5fVFjgKXROR+PVz0aA2LxZ2G3rYULgwRyUhl2MppvNqv
GQ3oZBwAoJLvPvCbUMeRA/0IBbP5F/5Z7U9lfgUmggZBAuhi+1RDJEI8lPHUh/Ot
X/Gmal6fkf7lDrTmwvLWHdc+iYO062BJVabHEzSrrsxlfADf4Bnwh8O+ApnFnpnK
8sJooU2LCa2ulvseoWhugNGNTYRsa7B+XH/F02X0Kmh5+HHpea0BHVwZsIBMCzAE
fPKw2ss74twlpBgO2D+mjABFfuq/x53nzQ1D1CQ05Ot5yuaKRnMKzyH1xmHIrIrq
YvMZQZjYgweGSYVX1ejnlU6SJqtrFFT9DCAmcj/nCs8Hx4ziIWReQGP80rXG69EC
kxiYe4t6wAosqianlmgXy0UIEzKVR5j15jvF5a4ipL5l+J4LjT9fyy0L41r+GZqj
AMBKT0L0/42bBQJjl923VhBkZWwWjuUyxYcIYtjWoOoEDMINSBVEUGdDswKXhx0S
GooH26ANAZSDWcBaXf5zQZwHJl5v5k/MIdVdHRMpH0E/37qFMgZ7UkBJqMrh8wIm
A1k1irX3/OJdEop6Vu8E9hr5Xj5UfD4ztt93qpKZavMQGSVBOOyBfxSqVjYOQVMu
lBqUdjNslQBfpfzJxWpQFsgpOlhmjXYXwpZwE7ijl0xWaz8sbgVpxQWIBraNkj1u
s/9JJQRsq3g3dfPu7lYJlaM/vJdPrFggenarhVyDYCsPaKD8d5dm/SLjCrnw9ANQ
2TAeeRbd3auK1Bp2rE1LX9N7uVQ3EBfN482R6mNvAipxftBjXNU7YjeB2xI1iEZi
LPB4mmNU3LC0xvieZrXTmY3OSHtf3pYzTusLyn4rVl8zs5ztRR/lxnYdGfN0x7JV
XX0EwepX/WFrpB1Y827TDV0m4AWFfQqe8/HFCk8m+3Na+si20hbfgnek/t57nXXU
p7Fhohm+mCH3KYtWHGXdtQIApS+7jqNVLeYwoDfb/CzutaHrD7Qzl3SjNVk02kw3
0FiuJqib/WPNiJLR3Y19E3MIQtOzLxfbHWEFzaeHVn4Cq0cKDNX/HxNCpYF+yJfV
/acdarTAfpq5SNP6ZtdhZQkREROrNXd0B/9YX5MSkWGu6UE9ORO89+sG7ftzBM8S
YPHHA9CyvbeZnttS+9IgyxRA0eZR0/ee+4FgthONsu9Uqlon+uU0ljYVeYGFgaQF
WnUTg2iFnwMX1+V7GWokCsqZEWY3crdb+VwnDn7Ri4Z6OvBY7UasTySd4qbtw4c1
5hj3W9jjvTdTJKerpJVft02B/CA+59RDwLTRrA4c44oimfzLCtn4EVmaZi3hVGYM
0rCUOLYrfs730jjQ1dNbWOcGGjlYqTQlq2Dl5FuBQFePE99hYZ2T6U1VqYoPE225
l6EZ+3jqTmrCdaeKTdENccJh8Zali6edb7nWk+sQXOWMrRQJ3qVYyfVcklZLGAKI
2xjjkNcH3t7OszZXAbr6ZcWxTFPMbfXWzvRd6OZyhoWzIr1ygk5m2yY3TwNAux6S
vpL9uKYcchNPyPdU0YEkiiDFW7xTq22UELJoAYU+hndIjfvf09GUH9rdgIKrMLx+
WygXrGBz/KE0ukYtgwA3CKm5uqIfbQ2iJnKuj6cE/TqnTM2OsxVgfE+rNzccMi5T
OaVOmc1bUX/5Dy5rhFKiA04C1SITc1vNXtzolHG37vvDNgFxFTOECL2Yr99UZOZr
t6NY/psE0pEYxdUzPGxn8zHcD6fXtFWLhYLuj1iQHBfLOpgzREFYHmhZj0M9XbWn
SvGNctZ/ArKbL8wy046dE+Yfy4vttbN7o58veXVxS2D8IvRflqPKHm20nefyTQdX
GagKeHVdDB/kCZBNZ8atZ2p4j5apDd+fLup5vyduqH93/oMLlgvqmzLOj3qNc+rW
NFWWDQWCZQ0xlIcYFYD9pt2YPFIIaeT4KRNXmJQTIHNpLcYa14EFyePaNE48d0vB
7gki461RCUujE5ck1YpONxeEXHY5Dc7TH+ZbClMZnDi7vCuCOLFavwZjpKqck0N9
Rr4HruCHFubkdPStwi+d3S7An1hm3KTWtQd9o87ZuXwkhXrlGB+ac+xOMpmypbT4
f8UPW7ZgaKkIWX30MweAuBjpPiP0GjC1FGkem3L3Bhfcgv31WnmC/2iAgD6x0UXD
bHehloya9XDyyGeaPRLwGGIp9dGrkPKtb/6eizFOWZO6p6sjxHkguR8Gyw2PQXX1
sPaoBgTVRsoDcLcu8dwcbqe9hIJBeKv0ShRPYF4QGAe8rrO/uSyX2SSAaMVn+6q3
npACjhQHpeD5mw1+lhZtUXy0D+vGPplQJdWwLZA9H/UAbmaAYo/YRWcPtmjTfa2v
JFwkLr5Spf4xyo7+QZaCYy8UaRY9MIKPd6O1JNUOqsIJsrbgYir/HtZ53Kop4akJ
NzWO3TPECJAxT16+TG9eyXF2uYNJMJe9KbzYNQmdpIphEO2WoDK4MkeRnbuy0lxX
ZhrFnBjDRiqN+5kOyi/5ngf2IUtBD+1hKuRj/+jmCbMVJoKeQbpVYuvgYojtop9m
8B0OXOhVq7u9ABrETOCdN1UZ0/z2Y0bWgD09eBMH27pRpu/Z+YBXaFQH6/sVKcYV
/IXvpR1pmGBGG5o4GaXI/s4AyQP6HKVK1cNQHjZ8jh/NQCwJCyNZF8CMDmzmgNzW
+cIOQ7yTbDSEv5/dhH0uIqjSh4Yy+w5cXSW+EPbWz7PPKEeP1EN5kxXhul5ZQ5jq
MB7tGOxDmmsyXT//BQQP+SpD7fNi1fJzzOFMzRUFuvgYCPHqRGZBcMRfLJ9if9Rb
wUUsDh2ery4hf+qpsaHPos78pzTRiS3/99tab9DmLxv04vb88Kvap5J13b6geGGR
KPbnz47F1w5ZdaN2TklZaTSIOTe1Jh+fyu94RsprJJphGBnsE3pxgeX4EXj0gjxM
CA6r5FjGuMCHddI4rqlQlVTUiBOoGG6yuDR9hGENbkQDAWlwX8nIvZAOcB6cOY+9
hYDbmZgR2k4JqJOT3EdqLgunE3glNBr7HoRl8YdxV+J1WorLWBHd5mGR+prGWqeX
URYgXTcwvESS9yLdMJISHvS+46kTYQPb1h4qSWsKQ2YnchZFXKY+U5JXFBeeZ6i9
48SeEm2YTY5mL2UJ4darYSK/7FhPplp79mG8bZ7MNB6ETuqtEhmsD7lB5Pl0mzIK
zUZNBsuibYhTEllNz8TLZ6lUheodSNcvCjQDaWIKeMIPwXL09peuB3OkeZRHNBlX
O4/g8mS35yaJg0vlgKQ7eVUqVdIfk9IiC++YWtlzT+PwFZetsyG/daCjNwr7K21p
VJ1yzfKtyffrhOtPM5+pZI44SVFB4+ycs2n9qtYBb3+tpw77Qi4jzZj3MYU6Rtdr
u0lcVG16OjICMKfHYB6DFuOVkrO6GW8yHvu4rBzpCN3wRmzghCdnywoIKsiVmZ2u
sYTLpwSM4SaVIeIJJqFnqlAPpFMNvtYGyGT8tY+zjJKQP3+pNhwE52kXohiLfG8e
yuevI22XSSPLHpVXYszZKTrmvrGkZ3qlsYVHEpba7/ktHL+L4kXs5Je5c0D89a/X
NzSi2rAifOXH7OFJOoGtm4ev8Sv3XIu6HsXfxlbkMFLOR04mvg51YPgX+j4WfcUY
vstFTe6lRGBijVCv5JMXAX3LHPs02NaIbElhW2vQkeVRZLf98v1qf+I+rrh2QYfk
vBM+lveZ7ys6IntBkdF4zvWqwJ36XhHQq1DZBoIDxvt1vTncDv/ctDVLLy3LUXXt
yIIuFEHco7Fmn1FNEgGr5BQKf4tm8b+CHgs8kF/j3a/MzBB/61zBydNVoYwRJlNv
CfYMaZqPU18zEJWequtwghq0lWc3SpnzBtdVdwY3/yoAZpYZ1tMawj1m7X6kSGkq
fhFOCSSRL18IS5ahbjErB1XK3RsoBUIAq1aFnKy5hnPhdTPJkdY8JV082DVIkHcJ
AWG3MzZpbY2GcLdhl+XXruVo86iwkk/pubQewQZK5lH4/Tt718KhiHEbIluWJ+X2
4Kec/GYdEIZokyPcRNN1hHts9wimUckm7PuGwSgFECLP4DqdImqYhFcdGY45sL+T
5S6eP27VmP4Hqz1cxW+Mwl4jVqDAN3ksGVSHKFef1KfjZRObxIS1rmGKQ4yF2ubP
8cwnP/1RrjvaZr2oglba9p6fvpl+1zRpPNNtzkrKIJ0GJCc3mawWa2V88zQk359w
dRywm/oeyIQQFvueUqD+deDBYjSX1nf9bjXWleN4d6ZmAvXY72iZEH9r6bc9H3T1
O+KV8YQ+G06GTRhx63uAV9GBgXWkAaTpqUGPRk8Pm+LBdAUfvDZSXxpBbSXeVEnK
Lr3ZW7vZBx6qo8CiG9bAqiTKd/brIFMukKUkXjv0Nsp58ruVia7bmN/WIv9UFR3e
hKKAC4ZJKKelJY7LSicwx4nzl1Au8rkIMg4JX0uN3fNNinI06xLahC8KEKklWdiP
Lh6AMIO+15gFkmhIIpIAUYq8r0P+tlCh49BiOsQt9f35gg44Go89Vi2CKPJ021eQ
Do8JHdavTLU/rfetCp+NtiZuTOfeFI7F7lAlCq9+gKoP7ei72rr4+k4Uu0MPdvWN
NoBp1eYgibWcD8brWVFmrRKhC8rrRugmyqf2ixzL5NMXOxobwHefwGW2NGgfDfoq
sz4zqYAcQdy1t69nZZk3xSCNtRkKAalk7QtCHz30JnoryuXhOtNhQ3pn1tu5k1o4
AZtPTGzAbkf1RGEr9oKjrbVnF+j9K9vzyEag0DkjR+tdh+hd8lORjDGuTfvslKxZ
HxcwmUWiDSfcK/g7rUGyS9tynaHMC6xiPWHaYjt7QWlWgNibVWBzKpSwPiAiJ3zK
0FMJjZeF5EZMRLipBRD0kzhM+Sttoh9JawCPrLnZhq4ZakaFZXSY901nLmM7tbzc
lM+Hg6RpLjUEGmC+uTmN1ajqrSrxpF63XiCoXRoZCogR9AXNFHvokUkby5m/fyED
CnnUjA30U3VWNAMEWGYA/jXV5sOgFJ0K85uxT9bqDY/O6QejOT2aDBAmoPTcglYx
TgR8fyq8ERXiSnjFDOLWJsol8XlUVvoSw1+d8Cn1SGCcfc8smUST/JmU6jigDCcK
z2va1ArzQbMP7mTGnIpZjyXnSX9dsfH3ne/cOs6JLEuowdHDJGIDhicPIaJs+e99
QMSfOxkZ8ZJ2xAoJ5sNCfGCrD5G1DcsLskIrq04QBS0gykgiiOBz4Nu1V/8lRjrC
yOW7/354vHoAp61rrHtG7C9s31fdY3LU/yZFQWnmVupMQYYC8SO5cqSW4RCGyJRq
fRa2HFqbp2RbcpAidXoyAVlb2CdU7eg5OEJaSFO/MCg0ZM6Qo4uTyukIr8beUeqo
6IoUHLsRP5uU+0213iuVZnN9lZYN2k6BpWpctf8e3c+QT0xT0Kw8LL2XnF+YWv9m
zxWpYsXaA4uKwMEE84e7PybLYqumuCy20k3EmID4Jv652j9g5X5ZIc3k+ksH61Jv
GhssOAlP5c0BNsm13AOx7eRlFL+FP9sNwllapHvy33gtmPxdmdLc+xsLmSsVIcdx
1qwp9eowSJGQ7kF3S1txkkPX+QEyxBJ7+qZlfSpCn83BASL0mEsYPLdSvraZZJTz
a3CYowJqGpwcPWaFRVp8p569DuaUxtDtEdv0Nt2Avd9SvSZGzztGSeja7dFUnk5v
8ygTVuiP7sGMfgzrZ/KBePZgVFvaNzhz/2nrFfN9XE7hNSXZ6+ybG9ayFIRnGiOM
TaoGtOL1Q9Opa0azdMlsHLQl/scm9ojKzlXTX5Wz/u36i4mCqZw3dVR50teK+Y6O
OJgHaka0jTecjDow1wKO701V2EMqc4NCV8ImkDAcQcQBaYv0cm2nK5J/f9JJlFqC
oDAxHDXk6jwFY3dFE78RV9dBVBbokjxYF6KrLPSZfgFt9IHwMHLBTEqNJtjh067M
TJEnmQ8bkSn+YIoLrT2yMYVEs0H+eY7vp7luMU6Db8vBpd1MMcCtgJsUrzA94XUE
KYoA3LQwYLxX9fCb4ggfsBz5htmoWjLCuU8gfNJb3id46/XrO4rAGjI5VFLDZSg2
4kEJAOz28F9HYL2cogmWAHjGFJXj/wnvdCtu28YmzPcelOpvx04QnwCssAVBzHhM
NGyEiQMALi6X8dNRw2frozxI/B39xIShuS0AviPbyJaVIwnFFH4l8PPpknn0EarZ
TnP/2tNyuW7m6Nit4oPFC9sqI+S9JDZlN8B0FyUbdBwYyto7P9Qv317i0ByZa7jB
q9gX4c3bliyvHzC+EPmIiWrzS/cyf4I9RlW6QjyolIj/YhypI7hOv4GEUv3cbErl
kKHQdey7qu30bAy78xZQFbifABY1AB5yduKir1rVm+IK9jhIOZDApzKK0jDhVy7m
v3AnyyD7lxLtqXMlQr/v7obk/S9iUxcByD6k+enCIgnLk+nD39tK3/SMxtGsLPxo
Y1SSSaqcGm6t1lOFbyEL19bStsEOsCiBRhikBhGfxIcZox7EDiAM9C1qiPx4NERO
k38VU2hptfFJDq+ITdo74uMF7+dXSTowkHhiP4t3boppKrqQ43Wln0KuRvuhFwnd
CTHpLJt3vLOWbSWbPxhnOC7fS8K/fQKbOzB2UKeA3BfcD29S+lo7iyjkBc1q5N0u
zwlj0b78KGiFX7Wo1bZk0Z8GTEJGdtVkR231uEasxueGVHEBPW18+ws6TtgAFDta
p+RicPOXjN6GLzo9oc7f25k87FYsDiCspbqDa5vnlQgZo3BdymRocu65Ld+z4z2q
k3C3MHl5El4bV+EhybRA9SfeNrQw/uGQ4KXm5yxItPyDwWi26UFlE/IB8nt1OodL
UbmxPIgP/5JKJ7923G4q+skVykf8ZJFDxgoQyDx7ACD1yJMAA+naZbHnmONSzyUR
G5tJKRSpdsRYq3nIzmDfBE15Qxuspq7sL29wx+JG3c8lz5lrKnL3Irmw53lewtF3
OKfPMYv2mK8tlD55bGaYLFAby6aolAas91SwUDVfciLIruRUYmzE33NCiDdwaKB/
CNohmIBAsvyRv+hDry2hZwd9UyWy2ncaSjM9u/ffZG2Bh1+dAiBu7EmzgWlZ3vZg
21D+3wVsL0vw21MZRyDDnumsQqtOKkYm++KstXXe4IlC/V5yuGhsQDdZq879y+dM
I1rKaQouRF4pqCl7m6tWugowBwcmkbdbA8/qvO/QiOM8DU7K1fhKWMvf76Xs7wca
2yfwHNn5z8OuZGGUrbmODLYIuTnYkmRmm9s0mbULjAd9N1vfnTNAzhwJG+J1kkwH
QxYNq/w1QedWEDz/+1nm0W7dZTio54tTkswqGp/x/28/ODBrml6pnOSQgrT5m52/
cns9H8/tauM0IVNvXI5tkxhBz7av+rhXNPMiKSMM6MOw0UIAtS3qjZvBbHPsM7DU
wLtgWpyfcBPrz34V+GnENrtE+UxCar+evmoPzT2HP6UMdsCiBYX6stdX2OXaa0yb
AB+HjnE4sQwBCZhuQuRgPa+2Wy6Na5QC2OWm1LpIlVOUHXvK6dfpnBb3znqilXzq

//pragma protect end_data_block
//pragma protect digest_block
hIDZp+krC8VzC/hbnWwR854R+Wo=
//pragma protect end_digest_block
//pragma protect end_protected
