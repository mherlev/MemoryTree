// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
qrCfBvNERF3S+Fxf8cirhXk8FEavGExHz3i75MlBp/wvTMF0cu1kX1p9dvQHsyyRW+n02GJt3BhX
S9MRaICOkpRBy/aMXB7yPou+pJAB1g0n0mVrAosj8Pp25/7Wu1DJR72qmPmVuPw/yLptCLBa6Qqf
CB8MtK6VXW9ERRbvyzOB3PQ+uwJoNKYIu7mUJMIUN57pMQH2DlIbNCUIAKUQG4to+csezwfXqMs2
qElP4CYfLbxEcioQ7FXf0EsQTvlPcKviyvobtfTajAPZV/67Mwge3GkFljjnd3gUb5DuFxiOnZsD
IWjBptL77r3f5RF+oazX7E7tvl1SDYr9Vop9yQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
x+KIom963aOWX59Thqh7MTK4SwdgXgcvKKtkFc9KfbkzQqW77MLN3lhqGAfcx9fUe+eoQWcwU3UO
AmCkOyUmePktfr8zr3QSHQNaOkk+u8XQEgwiowihvGE2XqJamLV6marq3CQGIj1p0tQS0kN1+uIH
0hpRXQjhZzaQYHEj0T66i73SnnPhtY4VJKcbGsRDq3Eg6Q2iMOcQZpQQrETQ/HBroSIeww55NWnP
7r6ulp8vJktCIDGLqGOtBTDNOOmhKwIN+qv3zX94yBxQ/Q9NvPeUqJQoukp+XAP5g+rq0tS1hMp0
NK13eaHfWZP11WIo62qE1sq7i5tCs24vMwrj20ZEpDjHwune34FQD9tVyN1iEJ/a0UyXQFL++gIg
r+kNMObKHoa5AzUvNfxILiOS2L4DV5fHGqDjB1TY9tVBbsNm4YCLiYb79cx2L1F6XPVmDW/1U9Ug
bsDQVbHSa2/16l2wBRYJK9wO1pMLAUA/3WwDozM3N5ZtQVdd07tPa7ACY7VFQOf+sA/lZThIVx61
PNkHb2Ts6xDk1bL5Yor8VUCLUMv//YIMftfkj26i4An5oi+fzi7OWbVxandUUOu3+dCbjPd7mkmv
B4EOF0mDHDQtgEkUarwtutu+GjhePSTDeyY46PIRsgpqm2tEb0RcIcw3N3tljFpJ4JOqYH4o+Ioc
vPRUmtdUsaRf8gxpweNh2Fjwb82xJj+5Yn0ax4Xpkry7O73B+AH0ObzwrOOHefii3n0eFA3bhsar
xunvdtOgKO4rA4qT2Ymg9qV+GOMWQOym6TvIvUPBWMf7gq0VK5r2jg+YYwoW8Srj0Fvnpl1BG5Aj
Kvu6epAhyoLYtLVIclpEGBiM/yWiIBU7W/SWi9LfXrHa0ThRAsVCtaiqBEc8bza1LvXAl3JaKTPe
iyRzKZ0RbfvHJzNPSax3Xn++oVkoCkb1va6pWYiyuXVon18OEs2ARDtNYkB70JPe0ZzwzTkedJym
uTVFL76XfziuEMkr8ngGLfwMbQGYu690VQhTHqpjrAxh8VDjuzQOF78gPCZV+kXd1TrDwVuTZwHZ
49+KzNbEm6ciH9GvgpBzq7Uc9bnn54lNS2lICJ8dBqf5SqeqqmgNIshegcwS5XiNwDO8bTZuScmH
HOXfuf4eRJImXlAxVHOf0wYP+sIrfFksjA4qe5ix5VX8CX+ulDBa88ZJHxCPLfWLFC5OLgN8hqyT
ksUuRilbVQluc6TwkIuvZKR7TGwS1iMI/JDgdl+7JfVO3Xo8w3dql4fGH2+ug6BOA8nLGCAjhIOk
73j134Sucx4dD1U8KszlvE5e+sYpicvrYZIEifXkUaNJMTRZyj7eAXobwlh7LhXWUJ1nIa/JG+Wl
rjZyLtFGohSQBzmWjm/JRduA8ooAFW4YFEtX6+t2Y6mKE9C4ia4sl76Gowqv1r2ONzOBQbbOSy48
LCnrIAChyGThS8zBEesIfKHPqoleRKjku5eAE6zVPW/rMxQwZtBNtG6Z4hybIDWAR9nDkJVY6Ua3
SjlUwWDZ7UAzyiOrfkvXa3TGSDI1FtK3iV/knlFOOBje0rnPFraJZrMgEUDNk7wPRKuwTpzR6v1H
OrHkRRIngshed908YZksUQT/zx1sB23ysfo9wD9BeLtVdMAR5Llr4miRIL7WPPW1h7PkQPecu+fq
nkynQy5RdeVi1C0Pi4+/VAR9eRTIQeEOIOb7xVFK2dXflh8RB+Fo9bpOR6FjU1x5ZIGCZvIAwAi9
Ch9VLcOMf/w9BwuhUf2uN4Tebbk0Qfk/j2pP0NGbiKXCquWB3sY71swJGdqoD+1aFgJ5DW54rKWL
oCDVdY55qHr6e0w1EFrB3wndg2DquU2FWwOKXoGE9rB2pc57x6ttg6UiHZTWYaca6OUzWOoFCWmr
DPVgLNUrnC1q87TY0LKwZIO7V9C9Cv7W+VBIKqK9Y4ngBKCO3VX0F74JdUlNE/BIIxyGhi41zI9K
n2dqXUrGLXMIEx4aVghvhZ8PScjDzL/XpqjWazB3xFEUvEbGDi2/agJcEN4YayA+I1nI44QKI1Sw
tShyu0iVdA613vcXoyUQ7Aszf1Vqw3uM9PbVFZU/QH+mrFA16VGuaTbcolXl1wiFFHmyhvpez1kD
1rEtF3ITMEsXupRZDgPM/WU9dQJTBN3eBJfdgGyHW3xRwYr2tU85iCuNbdCPaTUfvMpYB8eO2FN/
QI5ZGq+PHPjQXEw2Hq6IdmNelKR5uV5TVE9FQs/c63IuQS+Mc/OOwaz2woZnIYWZabVl3m5ITiNr
uJiNKdzlQGtHWzi9n8qylCKxVgrZbHLpYn7BeDPnNSSS/JSrrGoi66DXjoJWTUvNHxR1sO5CyjEe
zon28MDmnSUUOCnlSn8xbXc92ZC5nv/GyM+CVtVG5bcX11+GW0q12OZTBhvXW4MFbnXtV8toDmXD
U4wGzefUsARryxw7UwO/ApCSADIX2bf/7sRW4/CooK9NmvveG/qeDR82l6lCAYOsL1RChpEjzHA4
Jup1DS+uZ9uuFU9mvOdF1HM3uROayX/xmkOEKh119siIO9mwgr1qxQttb9sCT+A768o3A7xN6vM1
nqifS8F/l41TeyKUOWEGpjjim6PsKPHO2gW1YWBBmOEwuDfHG6XWR/xQBL2/QjdVvJ+6Hu8ZhL3P
0emyqv1Ff2M5PQaMURSoL+kTGcmp/YI9AQcl6FZ1BGDwrf2BlbTHkjZB3R21NC1n2VhfVg9O3ccT
1rLhmh8AyN9CdMyGt4xoKGDFJ9QW5hH2S2yl89QPHl6U6UuzwVQ0gX3Lt85rwgJxckyOwUxlKkhI
XLv7+gmtwrpcoENaYbsABJxdALczIjTAWksc9gz8sVmT4O4J4/AP5QBgQKxzdFkP/6JyhR5CQDA6
IT9pbWsj0yL+fHKor7TogWy8CWoKkpih4AP1fgQXq3SS1Olk7bu24dcbbxzffxOHGKbsbt2PD3H8
YSINIZEIBzFyzOcNTBGMbqGrPQ/cdJz0he452yA5/5V2Oso1QZEdXQzF1oF80H02eqSzfSfzLo3j
BCHZBPaXuVitv4Ky/k7vBXtYZbyB51zDsJkpulv/35dc3qmEmtl9vX+YmZC7Tdz8B0aOclIrHfFN
ZEIMcXJZXKZHYNU2c+tkKqkl5ypgZWCLoGrVcpM/L+vsbLVUsVq1hAcSu6OlCzA28z1yBtvOGcjC
vz+L+idFqbq1luDBbmwtUlXcrZ5yBZ+cRROQMDJ+6E32CKOYM0KiKDSbFw3cMQlhZZY+5TDypXNq
MnRgxazqNlvISJVymUIX3S3fPhCiBxG5HbDcugw5Q7whvP0zE7KWwLPsaWSCXaSzCQXKre0ax7+Q
XvEuGvaoh426iTkEjg0BijvYAomDiBUWWWrqSCIZgr9RimvIxXdQWPoL5ZZQa3FBTEC3UYwes2QY
eIZ+tk4LUGpeZOUTAL/Q16cP/Xrs7UPZyq/8C8g84y+h+5jcI/zRgeq8PCnTemhvouClSnWu0Ll+
iNzFgJpkgbCxEAu2BPd9JcQjz5wGLHAsjpINWfZ7+1YXZPZeizwEdIj01sCqbehtM7jb1aRF9CET
7PMCOk2lXWRtdx6R68wye2xPrbVVJmOnzZ6W31SMlrmwm8T2iC/gg/rQfE6Yulsxl9q1CTWobrFP
7gnHOQfSd8HEqoi1y/0f6BLKY974SviJKtgQhLNsDPpKdnylciHN5VrX4iXB0Y3Xq7OJanSyo4jj
kh0PRWuzbUlYXEdeRo02S9efFCpbadxCdVu63WgI3mYLuZJluDXax4ithW5kaaFlvd1wZ4Zc3crA
h0R8MKLYn5BbSBgN5RDHM5vq4NiHIBfN/o8W4LLoshlgejQxUGtCLX5IQNA1J+xFy5FHrjjKM6/C
WAQLV8btwWn8nIJEt6CpPj0orTtf2c7m/ioD2vloXD7MYuPf6KIs4zVjFG8YhAj/0/yQqZH0lQ8X
3tcqCDiACaI3rmb9/k0CJDI2horPjiPaJnMcr7IZ0VqC/+uu0CQnEtlCyI8WZuXuPVK0M7NIM/XE
GjARLmlNSXr2ufJgqp0x1WRlAfXmHMURJzN3AxvoBGTI8rJ8racrH4X2IIVPspTT/748NtsNAabg
fm4i4teIEwoDgedA33GrhVrCHjRWXuHHr5JliWzAYcMR5TG/hRv4D9DDKgY441UDKAk7gbmQC8p0
82A0M9q9vSvY2tgO2NAPpCBYN5/ym4AvGtcwjsE1MgvjVxkC7qJmO58KQnvtr1aF1fV4FaS1lEfH
bxNtoQCBpta+JxDQmKSN9O+sg3f63jGr4AeyDvLyJb+Hq60Qf+6RAGIeNLAY81PZM3+vNwAGTP13
AO8HWdn6CD55TX/B+6/iyXS4rUjoZqxWjvaI7aRYNaq5oYwdOByvmnAltZ+YQYpf8pjOFMu5Xg3f
6GfVMkxI4PwIoKN96HdCRpWEQDvdDzBMNIgWrddn5rs2Ina+lhGwcptD7abg/rsPNuMIrJ9znDk8
Y2ZOfNLFUQTIbDF0rFvCSnZdrAYI8FgTsnAV7/pcsrlr00xmuEfAG3wc5KaHiK5ly9rpHggaSqZI
ERWQVg5rJMoAC2Lrv+WayTo/oOrr4uxr0gX8yaZwd24kFt4FtAstBwKHNaFEoL7yNzKwZUvQOStU
IUlb7jk7SyAlpzfrL3KWMQCnIGmqo6QDALJXBS4w5wqo1lyavwrg5KTROlD8I600KVZwAH3GyegM
TyCmwRgq3GOTdnWCo8fLT3OAvq2FON2Wf/NOYxkclKWwTSQecw9OdnIh0Znddbu/kr0V84CDfADW
b9Rg8VWp5zdr+YIV261ehSJqgZBXjPNNO4l3HzOrmyzuVZrakIc2NWBf9xBs735MKqIFFZ9MNem1
BNMoGMc5Bpc5g0wR4EBsiyK7OVP1pVEN5aC27nE9D/tsvel2neU6Gk4qdkp3Nff1aCa6ONu1J+LY
p3L+l4QGRIz8LvitouYQ6LUKuFvbxp9NjQXW2g3hw+g6Gb4EgtYDk7Waq6df9srL8abe9nOziNLD
ITJ6HyvIXlyPTR3I7v146a/Ygty/4hhkUspyWADzmCV/LE0suz03c/RXzCCx1J1KFwwnkqm3CT4Y
QyeCMbg30dNFOybTvVdTTXq0FpckhahQP2xrCccRAjfJMRf80QbVqRqGwBXBw7UgT4NMVnfWhIKx
fg1eGu6E5ZEAJGpw0UZ4x592F2zkiKiomqk7uGCNNmPR1NxejwWMc6+By9A0MaIRgCdpgd0wk3Ju
yneJCCrvs3hQizLH2pmz4wELLbQuMXlsDyeIAjvvgenuE40bqEmnIMq99MVDv1lVoc5ub149QM90
+KwO9kieoSScMJnvLP76gutiCgmYdIFoMxKhwdHS+zIbknalIRAQ24wXq4Fx5MIiLCitKzzlka3h
+FnWdt3Nq5nQDmSVL6KvDPeOCtoBDhsRm1lwuL6WoR3YIol0pHGpm/YRJy7caKs720/nDT6eS4OX
qCmHrqhYkDuLwqrM/wyd8qMff6O1AId4HG57Bxpez51nk/FOmaqkD5l9nusipR9O5BU4VPcX6wxY
cHxXQGPgqoH6lb1qVN0U259lJ2iAPS2xuRc/P/KPclqQHkf8d9XamvJNZmIXNJkD7RKWFuWqCU1U
ddfHjmUIGErOHg/WBPnp+d/hLln80mQ14rI5RKDgUWQir8LhXZ7hWPgnbjrFI8XZwwDIu1/YeSnB
i3DvJKcr8/mjo+Ji3Eha0+T5SNOI2IP8aIjDwKizgZUeIkf/c8B/fTk1gkLn5tBdSAnbxptJ5RzY
wY9paL2QdpTqaOcvreCKJRRoWoQDulmk3GgZ0kI5b1qq4bPef7Q0bQGfPjqK/ZYfzb5XPC0Y6qWj
kILEtE9e/i7sjxRqsN5iSiCamBcsHaTdB88DCD0I1ZJKFPSxfmxxiCPsNLE8x2cxJphngq0aPEi3
INq5aa2ZqZxzme4yQMeDKfvuFzkbpAaVimuPTVh7ymYRVfVSQ29Obg9p3zvp4JCS2et10xiq0jS7
CvCp3pUWjrNgmpj23TGls0fs2GwTlX7FUq9ojWUfR+QDDc0oxFnB6aKjRX2aAT7FcTaLCs5g1n4s
UDOxTdg/xgejluS3vAD+Pl1WftBe4cTxI6GZIpli7cL73VGpeuQttY0VFtQzScxbLFEBnk9bQJEC
x2VjHKvLmSNkn6RNu7iebuxn62lB02pSGoYSFfCKhRKUPb5BViNn/pXTFp98ZcAshRyh0mmDE0fT
bEkLAcb/S5j4/+wCCOe6lbMzqZXUA9abo7wfqHSrnfxFbd3sPee8njHUhaoEPR02OpzvliuXXy0R
aX8TgllzMRiwI5b4+5KHbRppVoyVdlNDzb/bAPXdAqUpdubVAyGriNvzKiru3pWaZoFHk7mNocQT
+/CoxDP1uibWlLKzWPi4xxYZ5VAZcV7wzK3fUs2Jjt6ckWqwdrGQPS/BKBmtw+IZr/Xs0hD0Maw+
3C/503mc+Guk1BZQcxGbM2W/0ZrrEF9ILQfUaXjlYoIAcNdm69QVdFo7sjfPqDSjhpt8a/Aex6Ic
9a0nuSgr/4a1/IWBes7IwmLQf3QzKZDs4ZxBfn9TCzfw8PGI0RN6LYolVy2zOIXyyjaHhK13xYWt
OuTeTnYslDcUCJARDaCd3tOuEUkNJMe5qRAdT3y59zBmysytmgxob0+HfAUiiCcsiZLMU1eeSaAK
WVzbVy13k6bfHIFkKJS6MSiWi5NRJb7mtrOJLJfIRd5LfhDJnCkQlMLI26/sNiGtd9f5y0HPMfWo
RACyJjb9Vi35JLXPjec6B4u+zZUNiatlk1LmIVovi2/4/FXG0aRqnci0F0ahymscWfZ0RT1QEUoi
nT0mlKXltULyGWclPGVj1WhUkrtWkVgv517FSmH25rRhcEMIxHfVn3kgmmEVpLxikbI6eOmCf8bk
/BVQbziBEYHNuilbrVAvlUnk+uQ2+CfSmvBhMAEDMul7K/5xyi1eP1eiZCmz239Edtshbe4M4gDA
FuubVaNlBWppm8i4VxBU6PdK48TdMGWsvEzE3tbB5ApPH6d4Nh/lPzMY2IV95zpQ87K6YSfZLVe7
1ia8NAKcUSBCTDrc4FTC1VePc8WuzeNCMFnU
`pragma protect end_protected
