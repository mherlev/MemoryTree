// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:47 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
k9tLqcQd2vTnA6mjylOQFLnuR/P59TsMNkrW0hOxOj4IVZXpBTH0y3plF4KjugnP
44ZYnyT/DIjXo1UvCUA8WgMgYa62CGJUpEU6HKpSl/efUBoiD5zVDV3ikvYaK874
Ghj5l72o1ySfginriiEsvzHlBnFzXdHsG/ISCaAq8Nk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 20992)
dyA32HEJ64t+oUNlb77EDY4NQvY4hW3hvQ6KL1+CSWdRrpEzZTp6avHrMGYK0390
VLa7ybdRc1d9e0BxTYb3oailzwUyNcIsm64xhQl6wixhdcOGlBEofR2DcKKakDFC
lKVAvHctmM4MbRAXFbxNwbYMBviiR94axnQteGdbmj2N0r57jTAJLZKqBp/2w1vx
wPLdcjUM20XDQ6j42YHLPXBfdtq7vX88kFofR1QclvtdLVeU2ci9uFrAKruy1G6N
ZPaIQhLoBu8OnhthYEmLfOgEwjKbXCwOPwTTn+ALjTDPOI5/KrjuMNUG+IF76BMb
oA87cc3JGNiNYESDjS58lslWah1BCUZznArUT/G+s5JC87TUPpOzmh9rAhXGgvqF
qXE79OislP3cGVaoQygAB/Ho2hXkBZrkf0a+7eGDtF4nqU83vJFjkOMKqbAfZA1n
PRoEfQV74Rp5LuTrBrsq84Eo8hPcINOvanzbPeSRH77Sql2jp94OvJsy0RyguwdV
3aGkXtp+DIoY9nPovw4bgDzHYZwmwph66pU+Gu+TWDd43OwLylPutIy28M6XTs8E
U412MhXRN78/tjjAQknBjGrMY0dQaK4ecCty9zUiJsvyQ8Ov5pQTdKyvwdp4QxFH
kSfn2Ds1OUyS7HNnLihtqjx59DpTl5XpD6rr2o1pTQa2nXf0uQ3PQLYbNrcbH6MX
iRsfngtYJnaRXublqHzo26dV1qk9bvx4nrT70bIJZJEuXFFrVyxkY7t62+8WGUes
8yZrtl1HgnXY00nm3XpYKrY4dZ2PAi4z6K4Xqt+l6/PDeK6maPC/FepeFyrhOHio
uFxhUA3JjBA1bTfPRmWuvrdbZNhF52Js1B/pPqQc3Xj6r1gcbICOAw/w5T7VeuGW
kTDjplLfKasuLv3rrE6wi8u/j2USuDnj5g2bNiLfzixBtuH3aYeL67vLhdiC2uum
gC9qtOTm6lXKUsFwBaCWLb+2ovD0MY5gYwrRokNsbTF1Q2BAlVPABnLPmqBep/5O
PWfPtxrjS6+Uo7l0le2+hvQ6L4dUDIRo2txgp7+iLFt5FZ3m211iS5//UxHsxkiq
sjuNejax7+gcOnBWkQ2Dw6bBVV9HV0doeS4ar2A6GY86vLxV/YZEHodSaFlPenoJ
oZ1ktDBlnSkqru9Qyibt1yNCsATeX/pouZ7jtbE2IKoanowpVLAQCarX0Qz9lcUd
PeGg64iy2EhXvcXZjj1Yud703H1leKZtsa5H0xU3endVzQ7rFQ0SsomC0UiaWlCN
RrCdKg+D37WhP4ei1shNIDu9zyYwx+f0aYlH7b8xAFUEeRiA8exSweDD9uvCyY+J
FlpTnla2yZbwW8GYZjgTWTpXxA9aRY5EYVtnsvpkIeNmGxeFgbGz41bpvg2RrkAT
FIJoDkHFAnq8fHC88zIa7PbHfcwFS+sI6VQoArnX/6TdXLW3BA8HLw+grlwL15qs
2/BI1L8iOAZ0hDisXqU5q9RPuK6xROCtDLJjpbpdmH3mT747v+4nNtC7E3ztvrNX
RsmC8XUnEKjUqBRKVpOLwXhiOHJb/gXti/6HxRHYZOocC5sFPqB9PUcrq6X/r+Fr
Gbt9cYfCsYJTZFNCQv18Sto/zcolorvjxoDnBrvaTu8bMaRuxu6sA8YcOZWgNZ2b
hivx0T1fpliPL5XvyoBLciriTVJtuJQKqJtAsduphhdwPau4XCR2icVcDVBt/WO/
KmUXeO9qlZ0qVrPA7fKANpunDjITDU1vQpj0AFe++h2Y9dgj3vVd2Wc9Fl6Q6G6a
M+pqWl/Oo29u0kqFLndGwqjgk4LWmUqavvTdxvo2R764zdL1M+VgTv3p5+OXp5BP
egxcNiOKgutP5x+ZUnx8WpowHT7h0eZ0KcVIvy/+Z5Vt7LmFqaw5Ikj085oTG+9s
ShADeMksnJj/buB2FBNBgjWgSQpKlVOqzC8Un5t0zewAiBfEkzlc5jPIDg5I91rS
pk8TKzy4F/DsW6PWEKtf7IOV6WJeXd1n4/x0hTHxEp2VL4tOFq153J8ly7cJJkM6
87fCQcaYFZgf9yOKJIdpBgQaOdEe2cu9M1kJ9eAMpJl36JzwjedtVojcaeammo5W
ue5tZKu0WJJami5oyZ5trRmdBE0kAg7U0Tl0okPlEMTTabW/qSSGpfOc4fybSGs6
rlxmuoyEgModYtqlxAGhcv8ZODEP6bGbrfb9BUy76tzT8TWVwsdRvAqfeAxPfuxD
/FqRAEZWB5B2fu5+LgXwVjg9+23YAJXab+lezX5HBfy02VZ7KeL69b33xal0YqyJ
6Z93EqzjUOfgbgQx+Nh1fi7Iu/cTZKgNhKv232M/hXoSuCJ+CUdvLfqB++nPmszH
L6nsH5h279ThKTPTPEloS5hFD7hx1fasMxVPO+v+xbh3W3dLquOJ3kchTT2J4NoX
8Xsig0ZJYgr+xvzTYRVFEWDfwUYuQ8Vbf901mXpvxB/KEwcftPTeAdZ4Y7gYGOQX
OWipjHAHMlyAsj3y9EqvlhuSCa2h4sWosJzxhLe5ulVHVXrq3dOLqOljEwdnOFli
b6bhrdOB2CWOSLwn4AMINj2roc8NllECkh7krMlTAgiPOTMTnes8tbuaXwvqtaUs
5fsTeeGo+iOqa0v7EIlXPEm4Lbntm+8cfzUOm3cc/RoMO+JnGDn6lxfRpCsr2/Ul
SIEvCPda8B7spDLmm6DS4WF9XSL3LpySAwXOeiiEMMxK6INVHoNBZTyUoemcgF9Q
g/EIcCnbb2j1RJJsdFT0DhluOgY01r/Jdd7JxKJah5WNE/Mlg4eFvbCxm7w8PcTp
rTmXDXW8jDpKysuys2hkTFPvfn93uZ+PtBFiwBpTfgGtV1OfZJMpRWYYZaI+DvN4
UDk55HapZ7P7bVZmweBZKgVIRFLWa2QaQNMmChf1rLZ4kZgoh9t730a3bFBS4RJf
47PWAqH39Ptzd2vgcnPYytUEkoX7X4nm5qQrMai9pF8svOU63QNYgtNPLVsgi6VN
bs4aVYpp71VnIvKY0bn0IjsEUe3UZeCS4d3jWhRkPJWTE/tSojp34khCymJGU5Hd
6m/M63z6R/4hV/7LDRVpXGXB58ds+AawKjkaTaojDd976etAnd7SBNCoWUxfHrYY
Y8rzH3NSGY0GvDaLVn9yeQ4DTZL97WXvtEAXTzC3cVX/Frow2C4i3hvU/e6LsrEl
nzIYy21emyp9Wa4DUdG1Db+xsSSPHnrAQfbk+Igj5ZQ2XeqzrwACaYAwCnqQGGSi
Cw9Az+iRN6EiBmhIERPrOOxojkBrDVZ7zzrmrvlE8zldV+bqG0GXHk78fjgUnpDk
iUpa2Jq3oRZZlEg/AAsXgOPwJiCVKkl2eammyPwlZ9TJC4oKyr8iMGsvBu5hE7Nc
1cS7VqDJnbhRr4/x0oEZwKoLT7o2zJ4AiENEBKQUYfQVr4JlO3tSoL/lSSElN0UV
UAe5o0sN0b8K55XqgXbt88IDLc4ZedqHX94UNFze2vMLemYEjLR5IjMz2UhiLPWB
N/RR/c+wNVzbXtxUX9PVDZ3uFyZaknmiUvpMLATisAfyWc1Jcc2wOaCrk41ye6IA
7+Yzu25gt/BDPF/TnxUD7Zf7IpNhJ3gUtwt9yUcFLfA2saSj3v8o9IXgO3MnkSwp
dj4Ubak6QhCC5Y/BZPwmYm9QZFpsNAi4k6Svdv74mnB6la9ljoKmvh5ukRD7EQi6
rzThfXnJUrRH2N7sZwjTW8OUA1d72AfN/+aJcR0jmYZfG4lfUb3wpTPuFXKiWJHB
KDd9aHlSHj410ZoGokaVPK3vWew2DPkEI8tXhHfujZjvTlzbRIx2iuVjLOjZGC8j
sWtiu1/DJ+rgbeSC7baTi8lc1LMSZNZLMhCJUjT9REBQvYi1gmkVyZwyBYtzZhHi
tH5tolyIIiZIFqJmg5iA28DSPNnNZXxOGXEplubZjKMihPxmTLvaMz0zLgOtYqPI
2E8A8tz3XCCBSjZfiORgTUD11nCFyzaluILebWuHNG8LMDQlgBgrfu1qXufXJv6C
yXaRCQfA2CSW8aknYsboDwufcMioI/vSZ8qiX7+S4QX8jZSyesTQbuMenRMJf2E9
BhbKv32i/mihgGItgFlCMNskZkNwf3CoTod+YQcbKJZJNKAqHqr03U3Ikq96jJHU
OCJ6TYxpHaiEhh1tHmCI6T3/3ZgsTNM1J4rtRDOTf8FWTloHfTGJU1YVxxKQL2aS
at9r7FB5HV68cIgRWzZIrfgeKW/KAHaZoZHRR11ZTMC0amUyfvrnXttY2oCTUNAR
O4atV5lx3PjksgIT7wJO1iz5fxVYLqIRd79umtQlUsHGMVUt8nrO+DeH2lSP2bAc
gnD7LP4RFWXR1jJTWkxZz9FQ1RMrgVAx9ugtZRZVglN7Lk4jwZmO4tYEDRPwQ3eu
FMxHgMKUkPjvm0OUXHw++MrWh9prDBB5GtEUddL2V/LNKMKAiQ8/OSn4egZbgxbQ
8Oi0pAsIgYAxalW1hZYeT6kJ5zxONQvDErluyjiUqQTdh0NeYdpN2X5Clf0TfGk/
JcHSKmADrF91HQigULCTnOSR9+v3oLdDwu3Q8uWKZN7N76fiJEaLxjGLUWtl1tQ0
pGwayPbRJNxlAWvOibsVkS1G6ZGeLkz9zYwnt3c+dnywNPnto09u2YRhVp7t+6yT
e/tDq5tvAkiWVTsexlqS3Mzh8YI7L/EAd6vb5kW12vtvTJpeJc8TLBQdd7XUsxO6
Kr511ljLk0/c/SUl177LvIByMr3FFi2jSlxqKnMogR9VS4dsFOIuL8No4JbYliZG
c6KfndIcHjajkPeK4yzD+S2C9old8pE6fsWj7rvjj59FMcCX701Rgv8Bega1KPk7
P6U7oCoKUscflklSz+/YJlcUjjtyj43rNcVL/7UAANWLzvZESdzIwMapby0z90sx
xfUA+EjjIYKa9+CKLSEJ9HE0SqD8X8/j/sRz0o3AJMY4oAp8Ocv64PRw+qinY0Ii
+RHxc0t8c31GaqOeAlCJfoJmRxOo0vTHpZGxAibxW5TO4iCaLHD17FXv64THfz3P
PHBN9s/n3xGfefm08juJk/1q9cmKcfDV/lqPfhxOVurHNGCkAjcqU6sQTRfm2c+9
dXC0FJhjPy+keMSPKDHNE/0Kws2azLiWqvFgqtNAbHbmnHlRB8P3cs704IlQFJ0g
NuX5r4yiCPZrb56cYOOD5p6vPgqs18seiwcZDcKKjKW1jzkPrB+87gdevTfZD/pe
Xd08QSIxy98lqI8tsk0Sx2XIp11ilMe9KZtPKF+uZOEHeAr28sgcuUqeR2LVn7aI
/gpFVisU6SBRhwbMhXI1xvs2Ex5mXQpdIpmQZCBaXXnMDRP2fruyIdv/5rS5BNZj
6r9pfLb7+BIylLFaZ3264BQqLo90aQ16iwQ2bc8xzrAOzyUsDDfJeq8sg5BK19iB
smIRDg3ypYNJcsAwha8BNpc688p0IU9wu7QT8VCzpmxtAb1E/bg++/mtRM2ehC3O
PlSNBnrAwwSaAVY22ia183+uWg5fkR1BgkozHAJPGgRv6iH0K4QlrARg2AYIvEYv
7SOkLXmdlDE+C2scZy3B8cMRtKZCBw/JUkwtkN/0vb8oiPBZBiNModZmjMtTP3QG
K6c7PRxK2BzP/JfkRknWkBGiBCfJScbmtPy+YpYHItP3WtZrnUT6LDT2FdtURS+e
ceuJSm/E5Wz/kBcnELXYz1Nqf/XgXQXmnNwCq0WKub1YY9xBavyRRpKfdqhvNHdi
Ma+lEDLE1Lk0/bgAOKF/mxj6KnX+1whX8AJer+/irMKk2jQ6OTzOkL46WN6uzdGE
v59n1UMx6jJ2j7/3bzx5WisQ24HuZLGahgVcStd8Z0owoqIyTcIoIQftzN6CqJVC
TYKJBhCtsDiqGL7W5hy2yAbCSzL5BCWUv8nynw4vcKrHLp9nVwEgjUWzQogROcak
ZwoeZsvF+An8nGerS/UTegfT9hWeKx3ht3ePZH144iTehrJudjNGR9QYFC1Xh9bA
Gq1lvGNHDHCta48EIcUy9CZeNTAw5kC3PO64GEZn6x4uNRgeqiicKG1173C6hOzs
xQ841IRUGAfMi6bm9HsdLbNImb0Vu/9CvjNSBCX43JwnssKghQTd0deiEY/xB+8C
yXPYZc5t4/efgUmx24+aHjBLedF9/1xu2VCN7L2bjDSPXQynCSE+rTB3qCKPNin1
n91dKJI2LuLj+KHBWjy7D+Nh7EEB4jCdt2mdkbu2JcQZcFWaW7pOjhP8zZqJ38hK
CKNTFszayB0tZk/ROO4KWd1S9rQNqBqwL9vee273ZPoINTZ1tggxs6t2ulX0skV8
O0jm+rcqx4TyFbRyxJKV+Ti20KUTh8/8J9BupItlMjpXn+R77Fi8NroEtho+R8xC
HZEDeQs50M/Ipx0GmLMo3Bx7ai2BxbUVNTbL93ytcbjaHQfnJAkQkVvbxMi8yKLj
X/7k/613WvNr1AtV7gRi+nZ4smP2bZdewZZMKmdNyuwCn75TYWKt9SEp2OwXiM9+
eI0nbXSTSHB2uP5tR1H5FG5VGyfPtQ52NX0d3cq0kY44TMkvE1MYTLc+2tj2HH+d
sZ+l0YoLif4w4G03xqWnS5LKEVlhv+cdnZqkNyK6O0rD24IWJIv6SeaBWX/zi5h3
rx1VPwhx9eM4G4/T0KN9r5IxqPmdKY6X7CPo4N6xbZnEiZB79W5Q8JN+Rxl9slQX
DRta5MN5ryJoSZsawo35lvNlCIDM6iQAYlH6gIkBLKlSGt7SAafIiVoP0O02HfUy
Uw50ttzyRCfr2m/HU5/A04lJGteJzO40hckoWGx7U5GlzlU5SIpik85hnjUJm+IK
RUOyBDlzSILUs6vahGagf5vMw7Qfj3DoTcVasL4vOJsyYwzzerOV41dmYEyhnmja
iXf9OxyQ+N9xc3sEfWRmX28y73Qc/F8l0P8VDf5mnMtKN+b/sIuCejPIFPCA6z5j
uvBLLXcVdjrLy7iR+oGjt6Bl1BxrXSHDt3klWm7rMlgP7rTnzTa0tPsQWlN1onp1
n7yav9Wpko+D1d27BoJeEj6pYtSGYii6eSDg0AkAGfPw/ZYZYNTwtqShge1pnrT7
kLxTiTDm8nOodwclEqIEa9aY2DTTjoWLDm9YRYUDLanzrDHDKVZivu5URnk9BLWi
ucf49xQwqXiORDVVDIgeWcVUcfTfUFeFTcdI6KcsfA3tDoSeAmBQ+vTBpBkCnR2w
NnleFB1g37ModvS+obzYQn77cXK0Ov5ZonigNMf3HQftCqniWoDUMxj/gn4O4KnC
iyBWgQGuFFn5IRp2ODGdUPMyToyxTVlpEVjzuJ17Sr+wfk//wlEa5lcULFJdp2F4
WUItPbsHzRk0pKw8Ax9EVsXOU41x31bZkDW7WQzsg2X/vIp+I/ZfltHfKtwIn45O
+rtZc11J8j15sXcHfSY9xqTCisM39NF0JqeXODhmC2lCVp6i7XIqd4FLKdmJ/ywm
fkSySBetD3W1VB9bTud2YU+pA0hMzOc807ZTaPQ6fhiJFxcdZRDHj33d1eA2IpX5
b9cfQbSFJMhp4uEmGLwwhj4APngsVYAL8QdhF1ePWl4rZ6BuoazRtWdU5K4oEr4B
Eb6wR8LuFtftEcGFuvpyxddGFbmlitgxTQksrv4nrKznFd3F67dMtsgtOvDCsmJo
yPUKKLivzRND3Az5lCDaR7wqc2QnP7x1qr9dqF2+ln1FA1A0JYiVoYDeOzKaryZX
qEzVdneSnJ0Tf/GbnKX5eQ3iwzsKJFgCUFM10x061lQAXxEIP61JDEMYXmROIvYy
7P1i0q0tLQqSJ9nARMZujSIW/uCrPbNpWBs9A6qJMR550F0JpWsCpICBrxPF79hd
MHlMEFIUTB2g4Y6QRnJcyRDDkphYIUazFAO9keSRG6NxbdSNiDtTnrw7nzR5A0t9
bG0TyiB5nzdCjFC9AtEZRo1bpbTjlqNVtwNG8qrEVngC/8rKvs7B7dKRGjahiEQ/
2B6ovkD5wJsAEMLdPfJn+E4cOPjiNaBNqoWuFCAMufp5TlHVp8a+zm77AyblHeUk
60eKXqrXh0j1g5CyS30+YltObmu8Daot4gplrBGMNuVpRiSDD+ToekCjwgTB6mYZ
ulnc/jbFXzZjEacKEc6bxX5IoWCvDh2Qp7Byd8xgN6/3+Uz1YEbkZp+I0TpEufY1
7Ddz+91dg5e1yUc4J6LWfYDEVbsmGnuHoEaSb5uMSzsnazIcm/ig7eg2xBfyW1cu
yboO3hKWrGDRUIO0WbCV2wU6z7sT82lnAbSqvdI41e4iS1VeIjQ6dKuQ5Up64I8r
7RsjSjlkXsYq7BOs+N3AeRbUYj5MV/uCpnIsaiThUyMUBspmhJRFIPf11SqUWHgp
0OKoAlNItA5Iy3trGa6JoZWb/L9EYxl8D8dlcmcNFNxsIIUByQMh3JwTVWSDLEjC
+IdeojS3ysDvwnOImuf7Phc8hPiJXvoGzi3tqOI4pUJNcvBeqS1k9s5MXbYJuJ/y
RZJptvPfBYSVcsfm3bt6L4ZhGdqsNE1ChMTou845uba/AsVoKaOGLSUOhiDyBvBH
FCxofbGnr3nCwBET9JKIVoOo8uRUPE7tfIzwvF6vXYk40kt/93zEwg+QrIu7g1Bm
L4lctZMtwgyrmWC0cWJgRN7/cDp0w4wBgLkM0NjBtf4ePkg5gOpX+qpeJQvIde3p
GAL/eKAp9BoKIjjPSikWZETG1mWH1Yr5kmY7uS1UImOCP34Ih4hsOt3T/KFJzsAJ
JViKdm57VXFVXmwImPJ3dErdCceVP5z+NiEC6IsjRV+0Qo3Fnm5tbG1EjpmltlAb
mrBEzSVQ3MRl4vo9wVBF7yU4ozYrJmFpXBbl5WBVnkWYiFGgDO1hXsHb79iO0eNG
r4nF8T+HwB24MMzZ8zh3XMvG3vWNzSHEm7tFhiKha1MDPXb1Jfr69o7MP+kZCZsU
L7OmOytaG1/g2UaJOqcmysJXO2ywzA0J1jAz2EXA1jRGrzFhrL2kH/ZfEb3O6Osb
0URFwXh2rrmcfc//cJGUKHTt9eqg63d7T+qIGLWbNY6423BC0ojqwWqOtXsXdbok
lxm+sA7oU5HfpXun91jFCLFnoUZD/uP/nfXVfdQPuBt61AIRpF8dYSoyu6m3LHKU
RsS2p9rpWCgyGAooKVkEZiH9E9+HvGp0a+pU+WPimaswt9edLNSOOPUahCZlwu2N
SGjt8GQt+ZEcyPCDVLUIcswvYTBhcqTIgCdg3C2ETpOMFBRHsJ+fkWzj0YyOrjq0
ZDivBG4AdjCQULpnF7EUaFm/2cLuLivKyIhVzWuxpUDxgLHhyUXaZVYQPCGoYh2a
ZJYfV7cazCaNOvjp+7cvojH9COGw+YJZFOJ64GPSpRP6CiMCjfdF0VsUXl6vA8gm
JATzShLkhgF3CwBPXGM2xOAUEG3+iXlr7dKa2NVpJTawilqfFkuy1rZriatU0bRm
lUAtauD16iTdL7DFRLaBLz/y6NBTh8OKrlwr3PrAki3H0iNA19x6UvbtraN2BnLU
oe/hOru6Y6um9+r+mrf1+1+Rb2x4zaTRxinaKGomyu16QOWI5Bygp/vz3gE6NEXh
zfPsGTrJNMtGyAcspHeZ+i5Kt2ThEuwi9u7T4AL43yGThVbd2E5bmyFBoWsaHC7S
b/nfO/2EdDbrT9HHUudkVm+rnfx/fAiurx20XqkfmimLatnwiwgGxfx8P0CkRRDg
S8KOF2hARdbjGDGa8NZN0qB9YteTzy6phh3lW7D9rlj9eRWLJdxRHJl6PBsN2MEk
sA49fyvCXCgiJMuHdO6yAlOE9l8/k9qDACvV6tzOeOZf/0GWyKVnK74sBY5WLshV
CatqCutgTDOHmF1dupjrzFyIeTS7A738FjCkinAtXJm9YkBa5UljRzHzXLURBJJ8
23uxzERAv3I47iLQkr7QnrLV3iWunyuM4UzEm5Ngc3M9NX8/oAf1304DACbi+mey
23H56ZSdGpoJjjC2YdzQqPhigqwateMqIO2HmQSIpILQGtF7vEnnuIeUrXW2J/s9
c7Cap+/vfzOSuTLltCkctrXOMltgbmCRXpqh1+mXInCoxMvCEiaBywWl2e77dlKV
c/FgnEDGwP3oymZe07VkrdogvQZTtF2kJBCQ4jeiGIf9PbOgVQUH6yT+mOqwrBKQ
n1lytXzMjLskANS/KLiduFUEnIINUIGJ+Ef+TwcVGvpVXXCQeSU6JSr6gehkx8xj
yIl5uixxaslYyI2LKTQOb/9Uhp/c7lwuyi0PW7+PQa+10k37vSfUfSX7O2BO1p67
J91I3RUBDCamYIRaOI0kpzdMWywYp47VPFJoT2dBhbi/AdL/MP1UTUT3GcT3B+O+
qGXl8D0X1tnxFnTQGKWg0Yn6ghUS7pYsdHIVebgNqdoSPbZVdEXNatqC/Eog/iIt
Tj2zBU69odc7LJDwkITghiTY4WeowPvwU8fqQ+s6BWYMgXMiD0dV9Y0wYwd5QoBt
7fjYAsvet/01Llhthxt/XWOgolMbImKEYKYlwK/8xLXxFWYh9fDWzqrtOuDcAANi
cMFmehjpFPY3PwA/0Coy+Hz5oW5kPda93qVN8yhbpYx+zgZ9hPj7u+QTtRPOLQtp
Mq4m6VaZEtOzVn84MxoErfzOxtjnCxjQblxp6ut//eeZoXzXlpWuc0DUTgnNKyC5
lnKaFFxYVb4M49hYE8hzjcM+BmKgnFV2koS9A/znIN276bkECjos9Edq9TwdymGK
ajuUTEZnElIvf0ts1Df4wrirH2F8FYoDF3izS5dDF8Eb1Hjlwty1ACXALUvxYJA0
lHEuP8lzRWupjB1ccXxIBUFvA7OTXiAtdLJXDHXPtPARgFzF2x+4DZncN6jWeNQ9
u4kpMi1+A09rRcomFm38qIh4LZTKOSXDL0dh1PE+L7q6RRbnjBqD4iJVHphimZW5
VHT7MK+bIhD5bFohIt8qgbhE9fN+p8ezFnbaBFiP0A2eAYcem2CObeiiQbQtfR2c
tLryU+iSxJMGJNepA9ML2aWQ+ja8qPzSJuhptDEXwXTVj6Dp01pIcRsxaGQS71GL
+zLhb1yetelwKV1tkhu3hyYRYe1CNm2iVIVNqZZKOHqGZCceb7pI4XWXKT3E5o7/
Co4CvTsuzRwSHRZYhqsApT7LYBJsX2uqfnYKHpo5rx1G2PuR8VdZMEYVpXZ7Tiw4
0+g2IQI/KVfMAN4x0VKWk+FW+FOynLHAQiqxwWr+mEYNWnEFMnC5LYMm/1eaDEni
PVZsxCpBplThuSD8r55qmqpgQkM8mGFwhqNpgYCsLANWRkAYbjrpMEZr+8Df5vvo
b7Ehx9iedswXV85BBkvzfJmwCcw9CzPwleT2/9CDu7/Di4jB6n2cBSgVb4NlMkRt
JOFbFtcQKfK68WYfwPUIAbOB+r77ZH2L9qrv9rMX4IZEGDBz9AxSTtgr8WSdlL0M
lTmmEe1mDDnmW5q6B/aj7PW1ijEfc+l0K1DQmHB0Hr5j47tSMUvylWkeZts8zRxu
bnbqTmmTvpq/7wl6VlPGDwjE56ZuSPknVq1Hk0nfo6zNgwGdDwy09XmUbVwWkZNE
OCaYr6zgSk0kq+OpsXfmed75SOaiN2lYl9SR60/AFJZCleftLUNUyp2U8lvgLnP1
u2DEZrdPZBM6FRN9C78F7aTvhm+YQTuTgTCII6Osf9CZgsCNxrhoZWY1J1tB7SuP
vS1T2KHDUlFFw9o5GhynOBWiNkGN+fkSdjRyAiiilc74vUG+id8HsrG6+x/KJEwV
GmAFrN7YpkJ7rumSGesHXAHXTC/6fia7x0PNBTBREkxvhG0pwSuEhStbmz4B2/uq
xF4HFmbJfBkWA7SEkwpLxLgTh46WwJVqNPhjXLlRjRkaVQNSgCjYA7/ZxaKU4z4o
Zd1t9aE+c07ud1RwX+9dxZTLhqbah8lHVl296UvctnupnTSU3fPvX0s2XcWYDBD6
u+WEmjKMw5i8UcTM200y2jLHNMuuPipTrw4oZJpCkC3gd8w9awJ+CIxQcI8HWZlv
qU8XjdikDrTSjZ9YlHHM8gRNam4i4sIPxLUkmJVJCiRFmRbwgwVFAyrNkoEp5waQ
Naug91PB/t1nwKSnNFBKX2G4rnTNRoNhXbCDBVP/T0oUohL9yogOR6mRv0+omA5i
uOPQdbfev0lNHzDusi2PUZJoR2/HyfnREoNtmMnMaUm8iarFnkL9Oq2e049sPBV9
uPCgFwGe8J9zz5hhwlpAwqy/kSdRWrRtt1tAl+1DimgrpDTPjnZ6ygHO5qYE/lk+
PzRojFfFslaw1T7+MiqWkwXtMAKtOc6gsMHZo+Pt10YG5NOUKYWZ2GBl08Q2Bfth
j2ope5C+fuSSG8JVQjHpsVbPunJIuUiNylybkvwGDLSlat5//nFKA5Mx/m72Kuz0
MjU6e4FRui6BRiro+nb/53jTtEt8onnrUslHxM01BDFlJn8oROHT4ULmalugf+Mk
U0uXuym46ZCViJTDVox2o+OGLMZJhJzl565Dv1YsQSPrEetsNhAPa/wFg9NnE03C
x4nTLLPqnuwmhF9Y9zwyKXFv+VXKN01p02+soqTpPpLhM5ophNHfvbLICf4zfKvu
tJEDRu65XEgARV4jhet1sNPNIkn7+TQyXsaEH3rqmXygB1+5aMqhiIdn7TuuR0F4
RQ1VgDPzxM4zU3NbUb3ep1nSHrW5L29MYznRl8KnjOGpKt2o80GAdXXU7Lqg4wkZ
KrOcNEwLZ4NWk6pgB5XHNoEKTacMzj5mXp0cNMLO1z6NCbFweegK4+hU7YGoN9Rj
IHXL9C7g47suVfFNzAykaod23qXNsT3ZPPWjUk2tjidBx1y6HqsAM/U8f4lnZC1g
Q2Tr9naQhrVPNd4rnPDWgQVS/ybaAGFr89ibOQFxLqIhI35LVjmidDjWLw4CEx4T
QPHo1FJZFB3ShegUagRuRcevtssXd0r3KqxjSoMPTUBdSkw6lpVG/NxQNlXJuJ2q
OPOHg9iQLXI+sE7ja3d6ivkcTBunGFAMa7CcbmPkLmjX9Nm+JxlvfvEdHYHI9T2g
lQ6qaFZ9zR7bOEDW8+/W1o4xhFkKz+vmT2U0w37ILxBXzVSk9VX/A38Ld5YeXAaC
WzWrWAdZO7D77+cQpUB8Kzj1l4GT+ih5I2a+bsyzUUDxKcH6q77CMheeXBtfXzVA
+LVR1XUbj4adsY6T9RALcZP0c9ULT01wbw6mKsGPaJlL9ex4H9tIT9F0ZzmDDOMb
rNTtA71Wpfh0Qn+ElBhX3gQEHRNYLDWZ7RL3q2+B2olkUwpjyGF7KSvxvhWgXMd8
yMExnAGRPdbWHr/8EZAwu+QU/DCwtkqt07iJ1swjWuobM5RcfsZDOcsBkyj1et67
mK+1C/6gsJibIrOopT7rQq7aCTOa4G+Zu4AG1ZNTp2krEzdyzuxWFBU/Inpqef5/
IQW8X6WTrzR0vtYZiezeiIzqdXQbdN0P2cEWtS8HjqmEmR4HxjNggOhbpGKb4Z9M
B2uu/nP/xelprL2HMeXl44VHpLe2jsku7XINsr0tjsPqJ6j0iCWY5DIwWi7NN6Fb
bVFD4pSIPrPrAyqM57MYXsygTAv6uacE34g7KdvtYi2sq7OchqmhIrr3qNjIK4PX
FpXNvzO2cwEHNREyXEF2T+EBbqHqecLGDlPECox9whxSrBsgGLDhrL9GRpr5bR39
BG/I6vf+HIj+vAghKniImX1B9nLBTD3yXO9MCZWOS9APLLRx2CKr8kz7XZ+hZS9W
xWL0wn1d8omgadvQ6r8dcLuSPeyhxIq/ZDyeqGBUoQQYjvhyhOfqcUpSgV/f5WR3
Sy8GbrzwNDPeqiskiG9yuPqcmfg8SuQnDymN9B2wmadXxA/B5h3CdAnDoMu4qYLI
B/ivYK/Uctz5N88GyhjUcBtSCULrpMEHrQSdqanD014ZVR8QROwjT3mntdZBDU9o
YnGI2v5O3BHMphkZMFtLVC84/qGfh21amLHEfvSvN8EV6iggrVoMtP4Z9QHJoKAJ
QNUgIQh1IG1I0DN64SUez/ifNH0TjAQAZD3OJW0dKH6Jszd0skGgX0yV+jHcMWOS
9XqRIhgrjI0+JyPb0EyrUZZQVTBnPqobaSWw62zV9/iaFjNX4FY3mvLlA/AxGZw9
cS9b6DRx6RHtIeXV/g2QpQ59PgCV9EdGMa7SIpciPLykROW2EomX6uL2hCrY0ACg
2mMlsAZoX/S4FJ7d3g0n1y3q9b60rCXLDhdMOx8bR4sN9Baj+RWlMBxwTNut4iDK
XDOkpzxb617w8ebN8bjDK3nUxgdMw9M+OCx81yZa8d6Un5C/VLB5ACchIsLEZ+MI
bGU/vX6mQM1vdjjFPip8Ead03WfwVjzapMqCVgB9xjRr/BhpqpFLzleKgwbaiuBT
Hu6qqsegpaCMYTFdEBKqcQ7IoGCxO/ZVtgD7cqfh2/A5UY8VbVlJm6z2K3XqCZVz
TBT2ThgXexYbYPQcNnGgfRjFkB4l3WNyPNk+BlCCp+Vzn/fDE8M4bzcKgZLX3Wtb
+33On+6OO4Z/Ku5+yzkS9iKGGLSmHNGQCYLlEHIUhn7W5bEewjchc0F+ZC3mFeQV
5Ca2GCDERAXwVNEBvXLYb/zrOxn42a8EBSLM52lC4q4q2YihcpkRTYlTGEUpImpK
U8/04ITae0k/6Eg25/rk6khTK5UWSjzhpqA3Im9o4r4tTH6VBXWEE+5pwl6B1eQ0
BEDjlEureHPURDwKZe4TWUcE/uJxT1+q6lREXCqAMqr+N/KzonqRZriawIx/t60y
7iXBL5YpiSle/cbL0XfEvd17K/13ucd1BT1n4xZd+Qg6YPFtKH9pAm0dznGuv2FW
JTO+2eiYw7Nfr/dbVdnAJGGf2D59F4LtxudyI+Ig/0b1qsdeY73xmMiowbMz+Npl
2YR0VEkxLfmJN3E9JQ9GW5aCxayKgwILigKFqllXGz1PMTH68a2l7fUAJYP4ub//
PkCn1u8aXLcBUvRI4Iy0+N9qrf0TiEUf7d73qpBhQLDdozPLCpDk3wVG99sGw4QU
ugUKTSAYZyzX0k6pQUF5OIwoqkFVCNB+dxNzJm4Ga802SDTxmJH/Uks3MvI+Kf32
b/9mLirh8bkH9bVILvBc9vszndwRksU5P7htFGK22ZY4GXWpynz+jGsSxOOWfWX9
ZqfNnJIQsG2DBDK2nDjyU5SK3uBgpuP5gMQxKFjECKWH3hfgDfaBxG4ZTpxunW9v
7JPTeuoS2HKuNw60vvGXr7/c42Rn13Y/+e6dfwzSDpMksoH746xBBbMYxs8T3Vxf
MkzoHq4FFR1W5lkvmLNLmb7/QLv3RmE3RMpMiccJsA+VVd4ujf0p/YVAPamEnSTb
7RfyLo2lAjAY7kl7tfphNxOX0idLZB6qb4VyAg+yyI+t15kdHv1W6077VGY5HhoG
CrSmfZiTbNm9jJVMJara3vxs33rMs7m1whU5Vl4B5fbnFeVSmTUsntCs+2Py7Vz3
SpYVpCl5f08WbGMHm8O1a2Aeeh9ssOeUmK1Km3RewVnkPRfBmrmQw6hnzrCnFXMl
YmFrchZw9l/jWcEyszn231kJYIIE8gtu2lAIN+MftzhkwUiRzhQS8WN8TR6SU2lM
FL+e/f9YLrboWNbMXLEewcY4v0lcTnB4gwn/NpOzB+Nan81Sb5wZ99yaCzjOlFi2
9wqXGjN/oeyFVUg5PNwtdsv+vweVb8eL7MBuKJJZIDaQUwTl+I8YZ0Q3r+JgaO3G
+q82oXGWhCWeosrzZdI9rLFXVbqn5zM1C1q9R2/A284j3F2ismUT1Y7sQOwRIMwh
Xt82IXLYNZEJem/abKuyP6wX+QL6n/D3GahbXwb4DNV7gOj2TvckUlFgFz6k/r0g
dg1/2ayjoTwb0LgPTjgRc6WG7hoOv4aTllQziJd3yDYuWM0GZf0/QYiYkxuWgwFD
7FTIHl/8WB68evaPQ7a4xpjqyjU6FDlLtgPhoW187AChBRfG63k3QCUZMiPbbm2Q
GbB7LASInb6m6AY7kCvraZgFObB0aluIQa8mrHlKbBh3nkfwXYqvOtPQ0Zr8nhyL
cA1Rnci9J56P0Kdsh1DMvNjJ/BwaUoanNSvi/8W2SPYsvfA/ZOwocSK699VEnUoJ
edf8d7NwPzqPlTglq2n3tRA0ArEzvGsYOXivsKOaO2rrdtWc0E8K05RsedvcGwpx
0JgKbIwIAZ33NU8lHzZGCJ64YAEoXrcRuhf49015pmP/SIjSld+r/YTazbHJ3oI7
dfQUGmdYwkTjqLDPd0XVWnYTYUMrHC6Wk4OKOekSzx1AaRKe8f07KG7y3enyd73c
rLO/XEy9oK7hBeEgq7XWeCETw68FDKERJnTeYpVAPhTsYW3CWgfhmXefbVGpluG+
Sh3LPg7yzLrtuIJ2rPZIgkuR5ldm08Az+zjJvjTcExZEqdH3+S4G4j2TWo3GJN7s
7JknSoIZOsyPDvQdKqt97GgluDmnb6Jz5CYBXAIh83CyxdCI6MOO24/ny5WD4uvd
YxL45UjFUlZLhc5Ri0us4CrLIAgcI+TESRUzgtDb3LKcyPnKtlAuF/xKIJ+GuI3/
m/1/v8F1c/+TX0DGfRWThwPmaNEIHy26GCH2Wf232mRKWa1BWLOIeVH2wThtjKub
urVQfIy9u7aVSFHm4WfhMFjJCUlHK7P5gWruL6MGadC/am9D0cNMmqiddpEhud30
8nseKm0PvAfZzflfBn68KSvqBbodP9nDdwAD5kJqyEyjHtWlmxJxd2L1XG23oy2V
+W4CpRF3eOrfHNXSg7yjLpsK1L7eLk8mWPmGF2tmkfiOYW4UDd9JQHtg1E7q5qbQ
W9ET80QuOCZ3sRp8JKrFsTvRBe1UWkPlpkvXiw63orlg7PJmsq0hYz2fphoIr9g4
Jm5O4KL0UypKBpS7ikQyoFD7b5kHyFboCIasE92Cx4F8NrhUiB7rLcBw93qCV0J+
AOBj5LTEpf1wfk+Rp39MvVDvEPHuuQx4CsYVKLocnkz6Oe31bsbwOSFuuY1t5xnp
kF2jy2Klw9Y3/qZWNG/3t51cgG0bSQSAhAhBwhmkqghf/maDz2AepYXdcK+TysTc
bcCZGfaK6QqQ0310LbMw1AYP6VQ7FicHXxi+8OmCWnEsAU4BFEu8slPbEa9j/6ou
7UHc6H7jl6qO17hJxDymHh26xU5tcvVXPevk64LREsduGBBk+T2YqJOoUCL4rDMo
Sdn58tzoPu28iqa5iZ0QkNQYaaVlholl1xs7jvJOgKmtcbC4QKyHQGsNsRZ7Vl2q
IDlZ23MdrF1UqkGuvY8EdBcwMC3oD6ykYLlb4HdPOx5YXfPnNUWrWC/COlHHAeEM
VCYBg4Ti1c82Sc36AcM/wlDoBjwKioaPQUZUN+ClKjuSKvq/OoJaoGXcERp+N/Rm
ZGrcpdz257T525KlKfOot3n9x4yVYSzVpFh3bwoztaHsZ0rLhv2FNHBJJaJyNrOR
og19y25FM1rMDOSZ7damFAdlxHqab7Nd6flpVN5NVnBlwI5SSoUYB5VqS9rlNFtU
vii7GZsFGXgXFlB8AOP8F0DKgMmc5FM2y9qdAvrCoXxUByXzAowrsSWGR47y1Exo
9y5maKE+3LYLUnkSvhy4r2zIElH6ISpbXoEKaho+M5u+hXtln76kE36IvTdX/MKl
+RgVS8CGDEqCglOGFdq6GfLLC1FftS+/6gGr8svSJmw644+94r3tRk71GAr+hbe4
PtmVA1lC5Fp8PlDfnOyExVFhUFA7vmPpOcLsjo0YLLjGlSIqC3Pv/5wk8pxgsCEl
Ap2URwKCLYil0tuaZYCuozTkdhPDyMA6G2BknKaf8n/fPvi1d8AToD74wswyLmbo
H7XII+tKl0DTy8UF00flzlnD7ByNwz+FPvsenWDndaKv2nRpd+HvAbmhICk3ptLv
PE0Ui6CLguxI3gvoLTQahKsFHxiqslaIvs7ZdI+57zZ7nT3K9fA6YlV49xPujO35
SxV+t8neIV5dB77Q46BJISqF35rWAf3OUinjhd0pK0YgxKbm5N/nApbRAx/HzVam
NLClHvsDooLsFLOCWYVcGv67sDuKQFKwGM3CgWeJi1yxE4ZHFnR7sM8ClCt5yDWN
f4N5pYf4NkpxvHPJBcD1xJ3xNx/rnrLEzlzhaWaNbvpn+9J/yZph9CdCvCdLN8DJ
PEIsw7EqVcy3L7N0x4kNyQDMzHiwGZi3opBlUf01VwcN1JZREMO2ODE0U5+0ZHRH
Wqcpi2NWrNeAW/K8ciQVHl5/Lb3xjVn67Od8nxwYfRxeTKmXRyvn2FAGWMyth1bb
lr9djDZ+qNue11mObs0qbKusCNJznCC6PObrFydEKEjcyx+CBnp7t7QD1aNv53tW
lpyL1dFYOiZtprwhkhXcyzHb7C5Bzsj52NoQfAjoe8gBULMcxYo9c5NhlZ5lixYr
mim7FtgE1tawUiB2uJkQ/uHW3qWTVDiMhB3MOvBE0ZZc4PHAlNlAk2n9vsPSpY/M
9ea1bw6RDm2ZTeOs/2HJq7uiQFxfb8Rr/gajaQZ/e+8Omyvru9Zoy74nJJGXlp9j
tBIfJQ3zI+PLIjBdHoEocOCw2hcOqQeNFd9OyAfYzHK43X/xr0hFiGLrqFXPsCxI
OfmXh53m85rgAqzumABhCrGsCPTLOjpR040HArDHqgLLkH36thZYDJVSHlX7fTLz
xzrLCXVU72AWXK18WLzUEDUd/jgg16ocP2wDYylEOfF94+QQAL4wnZjpd+X5C5s0
BhJiJKBKCKd6X800iupy8ABkAX7ppTSR1J0Hi9xS0uiuyC74124HiyS8o3Nu+W2o
FbGpDGnyzHjVU38rL17u+1ebmLJesDjfOEGGsU5W+Kdd2q030V5LnWWsy6N3K1/j
Cm2z6cTjFTA8jlHuPM1IiI4dRVHw4crk/aTt1iGGh7wjHuyIRrsT5AiDY0+AQSwO
1yznuoZSJGe18Nq4qqm5+Nnv4Squ+2WuWwoRrcgI8AES058ioazC+rdW4+mW9RdX
S4W/q4MOzlEqdB/cVNOju3mz4oxJE31HW0o9YB3KuwoPnRcw3FFYTdfg3okNI9P4
YZAwdK4zwrHh4OpV1dzRsIupf04XR+kwNPvdw7K5/e38wzK7P92X6heZp1uitfme
SfRI14Z+QyUYFOaHyCwbrM1GYUyoOvphi09U/o9g5qBDhTZnTBvnJ5vo4Vy7x6LM
/bsXqvAGfDhGAdXNeSfic0nW+j4J3IzUxGNQj++4SpNZmuBbwaTBSU4/6IM/Y689
6SRHtEWWuOI1HKqtAq4r2nSYBkonmLHDp9t+hFqbcClnG3qFAoCJ2zEoORb2Uy3C
JQFXr9nJ+OLnNcdyu+jwmoMQKj2/0ik+ILLlhJ5sIgdFKV1YIl6Jgy/48SBridb8
0OYiTkIXr6jxss/173CoBKT3UYguligI9pCPrnSL+D0D4viKlBzlyDnhpBZScn9x
8bliJppisOvu9gquJ1rVOsH/CpTbCQW1HD2klDYQvx4Fg1vOSlZ5uUR/qvXVwueO
cG4DJo6OltQ0aXbkKbvWOoNzg5GHRQ0GS40y837TJF3RJirKXdJ0IPy5S6EeVTnm
KbY04IMj5TlPT+pYd7iA64P9zZta5mH7qb/o2RBsZxwjYS6FREe+EuehgkLr7B3i
Qb+jmMZnIddp+DtJWuIbNTrqcDb51/jF8k4Vf6JbOocsd8KGLmZhYT25P81RdeAW
pEpVfnF6ntokh6pjkTpLBqgQ4glAfjAhCN4ajxvwoynWuP30xFYDUBuObWItnJpb
YXRdP0rvH0N3q9IrBVdgpSerL7OVRUZUj1LE04WRvEBjpqH3OmhboaMj5qc9kvRh
tY1R9PxE4VdMI8zLLWpj3Lztn+Z9lTdG0QzN5qhJQZYQqcv9wFsCj0bSzt5OlHl1
yHjnwxwTzvk0eEHRefQ52TMYJm8jmrwIiLOQrNRbBvE4asVsBz1BwnAPwwnJG+Oy
FRkyr06Iutorurq8bTvQELf7OmdkXHQfzMl+keDGVtbLvTy40H4Dq8t4q53FJUv5
zxH2+Y+R3DTVpVixmFoAolCDOZIg9/jFKbNF5tBsNWDXNY2XHIrvIU+mzJ8Ouc8h
ZOdjN9t1mVxe6LvgT0arFbufJT2R2j6wyOYed2N99XLxc9GVwX5YZ1+fy5Eo/5QY
lJUSW84Oq83DaAUpgB19eMVxEZRKe6BWlGrsTgr2QBdO3clHQlhg7A3uW851Axvd
j2rd6Mlny8MIO/b4WYkhE/M3X5uYNR80vm3oC7g387vtrJc2bNsL8nSGL3+YF88P
v6OJ0uh3c0GqYLyamslu5WhluqY3LmipG98uWtEroOumriv43ebm5g5na2NoHAqb
k+QqS687XxB45Kj6nPEBXTYXkUokZewz/kqECmnxsWp+P/9Pq6VBss6HeL5oW8Vp
jdS66aAt5iDZge9W5nSJh/xMA1obLwxGTKhy1X2VENBKleCMhRh2DFPxiIZr5tBV
og6hLKkKiVvo6yH5Np3ZGKcO4Nm7bipS+wGSsuRYzZUV9JN5zyhWKegrXHS1eokO
YpqsoXPhTR7VDJwtzz/SWeVTvy4/6EA1LXZyUNiDnWcDQK0r0nJSBRdCSw/w49kJ
Ywxz3aE/aPBOoH78ISWgYxewJvI2ec2uV8s30hiCDFDPSvZqxhBCg5mzBWePGAW3
cfvhqOuPEdsnt3N08T/HZhWjXpb4PtbyFNuJbqay5+1aP5nfro5fEuET4sre9j6q
++Cjh4IGl5ax98hB8jLiS566r0ZyYx1h/uv41mvi/E7xq8tyK6q0cKbDwIGDQvzz
v4zeH5IDOO8aZpJARDXxlzw3fdP8pULyctMqIH7yqsn9VEAbERCPHLoPzoTA+hkw
AqxcmRcrHbxUbqpVSwpjsuyilDnBrCzJu8e+xihWqBx9QF8aVKidkVPxpIAdFDW2
l43kqvaicAfbVYi7kMaLF/ej2U7qKYnB8pXt+01uM+f03v0/ON4vXUhBMOX4Ygw0
2ECNmwZWQPNWXCSUizYIrDnsMqhqdYI9zS7c6JXLrYDxoxqyRHnH3o4founMCy5/
KDtbArA6UroE9a5ALp16k1N5PkdK40bgfQexUVctlIObaNjlLoBCy/15x+Mg+VVW
kDgBCKF7do2NafNLXTxcJvZ3g+q7d2GeUT57rDwNQT3MdAkumAQxaoiDDZJWtbFI
jIgeGwY2wETF8CrDeTcqE+gvhSp8Qbbl2mRXO8Eqm/Z3FWHmkLaKDiTtJPdfPp4E
W4yeW6AiZl4sbMmyuHfgSD1Wq+N1Htn/SZSgsOP8Fenx7VN+fJUai4UyhplH6rb1
y/R/3CEKmb5EUNeDqvvjMrwbwsaH5SbHdU422oh4q8fV4fDCXWJ+UBRDittGOGCg
WGOu+eGm9vHLSL4zlTrP6AxUVQTLDpM+W4IL4suCtAdNx3KB90byN/esyfpnGwLu
Ec3+Z3cCGbYEM1LE7bNm1zk4fxySjeLUYwwx5B2WwO0ewn9X42yf4RY2HRlOkKtQ
Iwh6pUFJRGTJXum1rYSp+dZ9FC6/92A9lRV5w3rtVp+ZRAfXKX4YxUatNZadZAgU
yrETXJ3AE0f5ZQbexT1T2HOnW+P+Gehv2s6slOYHuklOCGILKYgJMuKa6oD0yvpi
xOE4yIvJeYRn/Fsaqc/gyr8aI+MWt7eK/QrHw4mXMKu42kg5vpXMPH6z66rEL2SM
/FHWxtBw0ybkKowOWtZ+XmXTK0YLlyav1o4XI/4UYTZMFwAi7mn/Kn9aC2Qikf+t
MGkS0hYsH2RfangEa6sT8KkFlK5aZXEdS9mjAhOJioXTxPPCEpi2nhubluzBQZ/m
VVu0gjjVf30ZxE3z9k/CjD+kYai54uIfBAzEUWgGe2WvfJlgkXl+nqVtfmrwpED3
V2A+tfIerWrNRCGpXG5UoPtFBLTcDoq8vdN9w4xPUOBQOs7Xi7cJPbWZxKZzozVH
NcG9FbF1kSMq//N5EDRzDQOO7bXSvz0Mk+Ry7ihdPs2hH0mCXkwtO8nY9SFtYtzh
JjCwGSLqyu5YSwlqm28VsoeyIkRQ/R1zc46VyasmZ1zP/dZJ2/Rjc/CjNGzYEqB+
rvcQ7HsUmmOI+eSmjBTyXUjgPwoG6ighRntJSFMnfHwK/qwcBTUEO8dL9KyUGy5A
ywL2nIydvd5r+0BobYBvmGanl/hOBYb3bYhzsboigdetMkP3kCnNPnyY94o6sVJL
ycmWH1Okrr5HYFqRe9cLeuUvNfrY3fJNE4ZCC68GipRFZDYYerhSlFSIDf5ib67P
x9EQ0wIjCKnED/2BkHLIeNNUvg+FfnTes4QjW0l5hiIm7DD5czfQ5LUaMOLE7lbD
x/SqBc/41wgYzGGV9IL/dNn8yvFSC0fg/6hOYe9c+gsIx1aw1CriaVuDLumDFof5
PxStYSDAV+XfZTPhdYFMhyHvjAodFfCMoXhoo4dhHs/2fw/6l/DNCDwTBaGm4Zpo
LO/TbsF9VKMtiIH+B2y3lSLMpwbcJmrh2yhYTdqg34ZAppuSOf/OAupsReE5TFIr
v7Y8mRgiYPgXmh4wfHcvuKnIAtq1+nTkOl3HhQhPBGd0+/iTvz7SRbMsgvCE9jDx
ME/TjGkubU+IqK3LFsUuTq+w4LVvLiu3HIze2FWVUCEFPbDaMF0QQFFpfcIiMFWD
EVVuHefndpbBn/qmkHoDjM8EdDD76p6HXiNmWGSAC8hOg90ac+osG0xSwDsJRVHx
KqlmVRNba+od+QP0leVL6q0e+HzKvxnndUnB9c7W651COH6OV/lZpE2Whr8D+/Nk
Hw4s2w0UTOenrFOOXpvLrOhLlBSzhKTn5Qt7BUFUHz621xBe9RmEJveEIOSZfssh
tVaMethBb1Hv6F/N+m2bb8mRfEbI7IF9/pzMnO6I/9KSyJqd7w7dP12ebE+KFCJ7
cFIAVZd9TLInB1A5KeO8ABVUrKgIwegQoQ0797WYphHrg2CRphkRxdsUiYoM+aUP
pnTl89GzIwFHZgps3gr+mofyMCHvtTnWBJ42hpiYgTtIgSxBQTMrzVISAzNejjQ4
1nw3qX51R5iK2n8ByTTTHjWoFhWjeJT1Rpd+AGpiJBcFqBMBSSOHvK2wqFQ4JRzw
jwDiu0MJOFpprfIEBPJxiGkN7syLjVBgsZt0prPWY2jgfTFQuBQ9SfxgKWxu+pD7
iONAywkZ8kI0aMEbYFBgWMmzJ+rz4e2MQgroGpCO9F9qcHqhGcvN5J/ztMiLthfG
2cbNPoT8UQi16FmsaUJR0A+RE6bu3JZMX6nrFSJ/oJaStaQfYTEOoyPqJKW4On+F
SIwWnXkmOm7HLi6RSPgpO/stplN7gIS+Is/SNOqpY6PaSs6b+R9iaEFMzEWe/N/+
sWQ1MXNAxWT/LvGTZjf+Sc3Su3h+1+is5G7cMtxSgqFg/AEVaalqHUvLUAJQTdno
Ch5dZLwlBoVjN55ERvZump9y+qeQKZxnarMIassn/NtVtYXBPxBoTZdFr59UIpra
7zhp74hS3rEpgPQ/dHFDKWFk79p8a0cLdGm2jw94vabyCXRZPDuRltkcU8Wu5xBL
QbGFu7pT2kpl6jj92zDYw2rWlh6JCj7PPTN27ILMWKYPzXLQAk90Jee1cmK+BkI3
yNTBNIt6cvhzftEz6OovdAWb8ZCJrRKbJsRS1NBq28QxSSK7JLVJ1i/W/ESzn/dl
UJ4gdXx8o4SXYe5kxYGOCdqocxWQ4d/nZ8fzlmSBwJfJDam+kiupeP6UE7MuZAoV
nm7vblhzgQWgi2tnN2GNSzKoYu2ees1c6HyYL6Vzub95FhlIW4UNgmxsESV12BPN
8KTaWf8qvo0U7qLCzIqSzlW4mM19yCuK6FSYDDy83oYK1XebJ+l8wb9wikpZMgts
wXSR1izP8K7gYX5IMr9x3jKXxOJy+axcHGS/pMBTixLMsqfLuybdsQVO9L8BId8/
/aa9DoOhVn49Ueg9f5cuiMlfTP62EOLAc7S4PTR8P4+1HrAGyeWAW5yoxT7uy1Je
+lNsdemvrOtAbFRu4J2GcjBDSaW5pxaEupbD+A9Qcq/IjSBXl3kpLX/x0ba9ZQr8
aWfIqcZ+3jrlMJRQV2bYV6rWU7OFy/KKH4WPvdjzPJbkS5DWIWNG92CYUM/u4X27
vKLW3s/cr31usQx3UdRzxsVcViZjfOWxWwHznPN99Tg2lafl91NsBHKkHb0Y5NeG
opxo3Kxx2nbMiKyRAyEwLl3a13+0F8SHaTweYv/UZrbVauHQJmkC+gcDNk/RV45a
0WlgOmjISSEzmfetcwIS+tX8sJ+YkJLF547RFh07+gHA7hVITg8b/ebOurYEyoak
IbozzWETTqTkPoAG9wN7Qoj0OnKRlI0JoiUYwY1bIoqaUvwyOyxSua66PnhcZi+R
2l4jn62u87ecP3Lx5OuQGPeGNEEPlNumTp8buH7cdvQJ9H0qJng3HPO89nNn19Q2
uFydkKmZHlDU/X6yGgFRnzNKuwkx33XKV41nyDG/ZpoHj11PnRYwnHGBWIrtNNHx
KnCceoHoztRFtshr57SFeEEdKT2ammp24xTdhu6dkfyev4i/7inlktOWD6haA27+
/h+L6yt0P5GS/Nhv8qMYWRQokgNk7UaKA5WfhB9oi+Tr6Y5Wjwx7P0s0xPqZVAGR
boMKXvUkfkh1OWBRfyZxFaJTs8HEbAKwTyjTX1nA8M6OF121KIweZn1c5ZUh+IO1
3K57mPZCQxhWkEaP7XA0+h/QkiXvNU6Dj3unS1KBC7qQuqQVMRyNCeeIKCuxPea0
YzsUEzYfjll4MsN3rzn76zcxCwVy8zDv1bK+E/kFQRLnAXqxnIQAliXiRToTdfQ8
hOwd4thhKc2rPXmW2VxgsBnvnTIK2NmtLXjceGYs6johwZPuuhg+S5RVTCzrZ0yD
CLRKOyvF0QK7jR6Zcz3jqBkGU6EC+GUXMyrSChyjFqFHjG3ZfJdh98l7Bz2C7aX6
uuOgwgpaS/lKdGRh8oRQzaDlWnGJy9qwvHs2DgyFHkPdbZxjlAfFIQxRCn6I0CL7
WvsUkiyOtHz9JINB2iVkX7I2fgdoOH8kLcjPglGHBkr3uR1/8bhZGrvnHf0beYcJ
oGeMTWALP4Lwvvv9VtqdwGTXqAxdlMYWMOmBAVDFvDuePaOvI/bvq7GWxvNAn48k
mHsKHvc0Hw5YZa1Y2tK7gND/oMu2pV7lwUg2p5o1nMqtovK/CDyPOmMdT9KDbkGA
xMIWCzYnjMKGsNtl3aDym1Z3WuGEJ7eGHhooatxBNBmEnAKKwLJtZHdlxX3yYVgn
gXKd1qFbRTBXNYoPQGD0RxOr75PC0shsIIopgY18qIfbA7/cL/7LeJliSIchUX+J
o3K6Fk2AeDRYoy+t7NsoeKvHFaL05ae79qEqRzrUbABe+/ie2GJT7GlsP+HWXKLm
aM5Geg85J4qaLNgVC4Yk/hKP86BKzFx8s0UF+GbibQPZGwJ1Y1L2camCyPg4vXuz
H1SPYYrQ7cPA+o8UHSNISroGkr2VvZdw8b2VR8741MsZSVbAXjkKIRUzVSDcprYI
o4lm0h4zDye9cDPVuooXveCM9oJPLMehuWAtBhUdSo/YVeykJq0YMUOgUjD1u2PF
WcvpXuscxaC9ffP1Q1aJElmSDvEFbd/Hq3/rJf73VqNfzBjB/3RBKkNHTX2xP57q
OqQn1uL8OOG1hXo8pDEjvqQYXh+149yGVAvUfl1q/F41MxdHNWiJLsoJvZbi1UKd
QrZdVHCinUNv4eofTn0oY0tWb0kzWAbXz+d+2z6pQa28UtTPF0bRVjUogMl2QyX7
WPn1Fny/k4MKC2ZXQp/8cjDNi+v8ssFp6HC05XGHrSczSn6MQvQ5QEYrw+LZRJz5
0zTH5INKJcPOW6pmkujfL4xG4rHYCkFyKqUXG3vtqawtvfhiXx79iJc5c+4mA1sK
tXskvl+xuF+72tYpneWWDK270Q8vptZ/HhwCQC0N17lju1t6gkW9umSygl1n6reV
HPMYVanVRlnDrEM+GIXWYH4Mg+HzQOIfFL3z7SVi9ypeJhtGT4KRX2QDkj145wGH
8ukFtk4C6yh7XQ7H4o9VALMBU9kbTkye7YNBuyjI9VQvIo0z1noQUsRbf9Msu+h1
BFFWVRNeGaGH4KUCc7V/b4hWFKuQP1pd9XNY2TfI2Ca0P3L3oIDOjLCENiI55+H2
DIsKfj5kRlQPR6sT6ehNeQihfJiDWrji68Deselwr2BbbraPwP+K1sjlGHZG6abg
YVDHAb9FzxmyLMFlGHSrP9HhpjwP1Ri3mGiGaRMeegZIkynC5Vt0HXzg5r9N30gz
GevkYXfMM0P1tQamCMjWYpSxflTUQGB+UtP4gtVfVBHYQwrCf/v/I8I8DpfaTOBK
BtEXub7N2P3zuoj3XNnn56mAGKRh2hI2u2nWWZGPao6bMkFLGj4P9EdeWd9HFM1X
2/N6UnSNzsSOeqTU6vYHJit3YiWvuiE6q4F0Ohg15u7HjzTN8NfWshLVEPlaw0Mc
bvK55caclOt3ccfnGJTfoLm0cMjVXNA+rfXrzTDyJfMZ5ftpRY20dcRd82DRZ6x6
IiYDPYUb8fMYh4XEGqKTGc/1isldJdltxsHsc08KQ7wEJyu4bNir0dqdnb11y9xG
uzXEwHHKHzOmSaIooicz89U9rP8AK6ZeAO7M9LiAwVeQS/kyoYsfcJsMj3MHquxu
OAsXtW1cKBvMcVw926V9X+12Gl3YsPa9Tw4KrX+O5iJUO+GJRts8RZrLkXTlnxoe
7ggXZBKlZ8abmjRySCDuid2+O7wQonYxIfzEv0OMyBDga9K6hBz/wzLG8BvGCrN5
OXaDyZMu7F+KvXbvM9fAEQ4vBbuvG9488b9djcgBuWCvA9SodDRZKsxZ+I6esBtr
0GQQh/TuFhSBJVA8eL/IP1YfRyKB8ZZzyixy47BSMp0sKKuFNs74mQfT0nZjqAeB
ya3GtKU4ULTaops56c6marnySqwb8YaCHYTHJBCypsUvr7UOFpWNlLHB96zxRREk
oR/CK/cz2sqLDGwpv4b1DbJ5iNCzA7G7m6cJx0g6EKr7jZf2gllcU4WRwh+lgrgj
oC+EiYnyMzXLDP1ExUIg+MIFNZuxFE8Z2FXY3KbjwMEKlfwVl0MlqcHM8Lh/FEWP
UVLL82qFxR+mmBe4wZ+9/4HWuJjIjoR6ezqf340HuN3ttkJ9xm1dxEcvY9j45ws7
j9LwcxeyrzVqcJjN76GQCgJunQHyEKasW0MoAighjRbLVMz/xZnBvMP786q89/op
gVrYwVnec49zZkEPMh8gXbr43iE24sDGgJIw6oCsAWCa5MWqWSIwq1UDSaBlkLWf
Df6FnjHGfjQ7mLP6EmTJHGSuKlsCR1Vf2r2S0bIpgSmygrhUOtcHFOM/T/cKoK3j
/dAgAqWP7x5n/DJNg582wru6sWBNpMmSJZkajsFP2xe4EiAuemJSacvT4Paoc2+T
2GMGlm30l+UkRcbaXlSEdWE6L/kL23wI6Y0UTRvPnf0XVeZOey7aViEIAcCGAx8T
wuf+x4rM5p9Rz69b+3O/X5q1DgNxkXlSGiBvAIFdPsD9ynEplWDUP37kR4kllAn/
pCM9uGCaz03xBjByy+3EIsDkzrYvzD6Jn9mPnsQB7zaI25CITfbghKUimFBz1GRw
P8/mn0p51dx+9xWfVO8klnRhPmYf+hIhJE43kVS3AQLpMGoNO3LJhwv4cRaW26+I
4JSMH9R0SKNZ7FSl+HhJjzfn0CbQWJR43pOt1L9aWBDeKv+xmMJ3vZPyY2ZXgW18
JQlHGR/iL529zXkSdGR3h203anwvDEHXzaOrgDSNTH49t1f6Zzl3l/3xOpLde1G9
GLbmIRNc2IXQdy2/1zFnhQwl5lKQgaUCQ/F4dwRxtif8FOI7FmgATj3oDna29ge/
T62goSfw5wHVY/mgyh5cR71H/CQXrOx3OCVr8kxF96uuCT0NVOLL21HQfR2OcUrW
tBwfFxQo10CU++n7i+eg5w==
`pragma protect end_protected
