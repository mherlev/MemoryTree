// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:50 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Cw8iVGtMzjUgne8gaLjve3k1NdwNekXjZLc1pB+Ols8O9AnRaOhMOqG0I+rQmL/W
sF5AZiQtluHFE5b1SEUJNBkUEnIuiE8PAn6BnJOCOsCLRqANuc9hs7XcrrOU6iuE
4GSX04XXdvPMlwQ79UKq/VCjdK7W3MJwhq9WaYtJQi4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 27168)
evzQCiDk9akGB3j5zPZsjgVyhGUjjBQs+/vlW40iZGOpi8MJ+0tWOgjVxOSjC1bd
Q/dEMwf337ePL4FbMHqZ7PVOhjRkrnyiuU7cnfQI6VDr4qxpgZvKluW/fvQXZYlt
9K1vfMijH054ec/Arak7ahU1kocPAm1k9v0RcEF71W5Q//v3U8DvCrTUx3KhJcvP
fLreVz06zIaxGv5a3YGSL05XghbvNNAg8eYcP/3a8ge+TKAzryJpV2mxyNo/3xwA
bE81tPQcVGwoCiRCRww7iFkpBa0d5eDbUmXjk4Ksl8YG2mhzzB4/3JOmno97RkM/
+6RqpZat2N25ClyID1Mp9YgeRSaSvxEjBUMu+u/6ALz8GU65xlZpZV7NSLR50RsB
i9ueTkNH4BIUF+cZXciIylm5yRWRg05gJ8L/t47/HYKkOWFi1alGeJDsKDHwYUc2
TCP25p8DMkTBdcMYyb1GVX+Hm2dmw04bGCL4mFSKg2+f/tTPNl7bQmxU18DXx6Y9
dWUuukWcZkrwnLPnjoGxM31FwrHG1xzOZMY3Xq0NzqjFKTSJFMyZ+M4O8Knz2deY
CM/OJJ7wFkO5CscN9Tec6ckoGsf+ss0h0J6MXmVYPdd7IgDbvfUe7RZby8ju/9my
t1QQHU++61BfFwxo4qJfRXbldvLUOjTZeQfpK/MphuRlMMINQLBfOXISWrKbC3vS
sZMD9gGrljh2j6c9HpMVCk/H+Yqs4OR03BOSx8Afuoj0TKlacWnGsOelFwHwOP+2
Ljim6Wrchp+FOAVIcooyhqV5q4PXvKWIYL8gZMyBJwgZAAPAnIHjEASPYvw49NPd
jENyYGPYHb1abx1McLB+zuhRZ3/S1uU7GkT04JsaMJWyH7602pngw5bnK4NbzqFt
lr4E4TYwdAHnZCKJ/b475gtAbxDJewlkQgxlRj6daNaojoGkQfjgQnUsoRwo7V0r
zDZTBYxnER+FUr71K4AvgTWvt59+KaKgdoXiGmAO9vAWEG+FF+MhIQdyEQ6rNjRV
7nJX8/bD9QGd++JGL1A+cMDgkJrlT+dX7HSrmb0/yEfkVxqgy0gUMhVpPPx6rA+3
Dhgw1Flw8tO4gCUqvzNGaP3LwJD30MgaV3LEBDSK0UJLtgT3kC73HRpCOByE1J1o
bML9Odqvo77mzVlZ3BcbxRPfvJITOUZS6e4MAEXkECzA8lI1omhTEJPnUSQmM+ww
HUxLw609Ac+o7SsvlBUMXX70McPHdXdaJvGGwPTrwOJTjwIzs0tVuHfWRhE2Yxnu
GnEM0Pg7poe011PA9qXaAYa+PET53kZhQNTkOyqsDT4urfiGRgjEHnIgnqrmmCLg
QUmxpXiPlWFkmzphIJmKvtrSCasE5Teo2kSFYAUU0Lje5eIntvd3V0q2ZJqFPaNF
IMqTv9fMMB74NTTe8Xb0VwqvnHGdVhZga8B2EX1UoB8rwKxak109+g0YbnxM37hm
qUxcACAdA4KMKOkt1zziFVCq/uvjEBnuzsmkI0HU+rEEmu4862eJ5JmEybSb9x3I
NhTwz+AOc3S35y2wR0n1EIozy35X9Rn2AXdDrZMrvuxnxbV4VPa9YfFXZTZOS+sw
EYXWB8vF0O2k0d8Gqfh9LLy6N0iljEiJRHDOSkJxaATWaQzLkTratngV/+ovtGt+
/fQp1sBOP1d+6eIRVnLn3JLxwAFXFTl9Ma7tGB5fCv6t74o4ZijlqpMRHgqWyEBJ
l/hHDa7AeChTUkxK49JVtpZ3nL2La4z2pYTKaytjd8SOEYY6PGns9uVDdJkLs/cd
mzFJyrV+FKHdap8P0ZJbzpAr1nJS4GJ8yxMgUGntjjZ5k+DMrIk7oDJ6gF6RG22f
Lr+cB6XPtZnESKEOYSsbvOjinGCuyXyOmPh2snVLLEUEPOjdVCMMz6mBFjqp9MGG
c0nf3wQDTnDscFH0092eZaPYjwjhv+1HSNfDm89z9eTUyNgp5M3gmlrZA3CQ5W21
ulzwVH02GtuXExLtv+SvoVXyd4DvDdWE4I80l+Vo3Qf4o5ygA5/uWgoKjm7xjX8Q
w7N2g+geZBT0c62uYvsbwVBHkOkReIYfcQoq8UGdLaFzVB6TetR4p6qIQ0pqSHGy
sLHTVpvLNv8yIWf78GFZtQkED68Vrf1VIYnDE0w7CfUV5GZ7IRSzqLLOOgluO/uo
rEpI7zKCO3rKaX3RhVyJfnmZYTv6x5TiG99V78vLLH+7KJVqEB0KVgGqpwR0/5oH
uKSVbTsZO97VW6EW/qS85PVNpwRZpIXxS3auJNSf/GlScfXGBYIyGae2wZib+Ps8
UWvX+bv0c9UYSYynrP40w+CGZf9Y6BE3VXN6LJB/SQ+SWaapyyV3SYpjZ1NfLfH8
RwzEK34b7bojyYnSndJCsfspIllktB5koA84yMjK1d55N6Pj2CI5APEj8rj5biGI
rhpKyhvLL08HHI568oYofBWg3YQKSWw6oCvVCdp5Rlb/RT5ofvy+a6j4eonMdUTz
XSMBMgNm25b1fTOFZNjEoLv5TCGXcYb1v0HAoL7XXx5vXYrtehF4u+cUipf1RBdq
VjjJ95yURcUYNjwxwNQUr2NVPTFekBLGulIaWaNFxiXEtDqtBQ7/LnWCmC+kHpLa
sbHsvj8Adlhy+ljvIjR2SG6Y5yJxqmDrlvZ4pAUYWCZm5myxbhhcl2pmmppzJjRy
3H8QryvKN1idNzN1WAQW9h2NRmFEmzeGM7GvUSz5/rq4aZPmuHhcPym/I48SmcJI
rDsuIOqoQYO8WPlIh5DX0LzbTxsTuII8jJDYxgOpELpJb1O9WHTS7pLDbL7fFvov
LKOJLhpRUBfYeoTt/QW4CZCH3JqFLP+OJg9lXymXxQiSoqX9FiaJ7b24hImT9iXO
fuSfnp+GhbUWjpu/GCw6moWv2nkglNAPcqeh4h1EvxFRwXTXlNffwmZKqlYaLkto
kEpJnEEo/3JRZkRyWgbr/z/WG8GmjNMSKYrp07gZXAqOAB+B040rZ8lrsOKXMrDk
vvm2Wyjulzo/IrPwhqhjlUodjxVM9+rua9KTPFfUDZ2771vZnF9TJdc2DgHM9s1E
L92y5E4iOl864AXWw5CHRX3LSilXzy0zxIXk5gnK7lZTuwmIYeyB5/6M1yrwPpOx
ht+mK2earLNW5NFortusRXrwJe/vJxn/eNxRjBKyrlaujtELNNYIxKKRnOdJV211
oxMmMXdmViCUD6Sck88KscrrOFDVzp1MofeiSxWmoeK4rhYWcDVQAtuQumPgsifO
MAwqNnSvPzEj6lRFJPRV75/Xrs58b7jLkBKe2gMJfzUPvnvAxtElxla0bKEumWfi
Gk5i5MDsyn+JS/OBYm3pWHqtegEqNwtImBzKDy/S501UKsCKUK7PvN0ATxMrRr9F
hewuXEXuRPmQr+nqgT9ruRJ4nR1yEh0n75M/bYNGaY4ZNK8OmGuYAhzIqZkkkxUh
9uL2djgk5LhUEsQKp5VgKS/zl03n38ddCMxi/B/gEW9cikjR2CC9mgUrKIVsec/z
cAo/BYI5kxEbGrrOUZyXEnvax5W63XTWqTmodlcFkfrZPGVFXV2t81IYVgxxOOgm
7cKheaT82LfsXi86E8vWSWdEL0ltvp0bnFz0MJLFCv9+p6G2O8aGsAm0QxgSC2DL
rFfxtTcjr9GHngW56hs/wN37hmMlq/M5pBVrGNAlWgVA7/L+ux3xvAlZFuy4jpUg
gfBVfT3CEZ8Y1j15NJ7MLwtHts1YMrwhGbBdtsZalvJy+WyvwV7qPeh4S13scHgG
g525LuV1dukWTnj/T/UFJePeRwfZ3uExfRnrzkNTPvr7Ga5ArErOFuGdeunT6Aib
yljutSN9rUqI4jXupuGD0IuNn2g+Z14QXjOJTyzEwlrICD8TitwFjNSBaSbErZBx
d941EMIrgitWj4WKVHqursXmqNFskv9DWGdeK5CFPn6StrYdDrsujOgesYsSSVtT
lDfZm0xZ8bC+OUn4Im79DTBxkdJXm1Gaa2GjnPpo8I6xzG0feOiX/qdMAw3zomCF
w0T9azKm1bps97oxwoO73fTaH9lVKVGmHaMFfctsebQySjsvrol0b3ggH3MYOZ6N
40+ZGzTtwkW9LCfZNJNY7qbwIGj6XYLdc3izje8oUP7+3bGmkd6BJyYzG13YJd60
RC29lPdI1dq2gIiX0RD2XsKFjt4LUHnDEKv9r9NT0uhutq9MuLgu3bSKX0ZaWV5X
kRWnoXWRxVmfX2OzLhGZJaM/RaNjEgrxpyDcPE29xM/n/GKBOfGkj8EbMKLB5WE/
0kdjxoG6DkL370WpsCMa4h70+nYpFuQw28rhxlpS+9cse/A5jLF2u/HLviLOki/0
ZX4+7RDc6cdlGimvy+6hsxkhrE9Xz68vUUAIEiEhKJyuzm6HtgW8R2y7jmZ4d64/
YVcycqW/AlUPOAo1AGteU6mzBUTZLA7nxEzRtv1GuyFRlkNzpZ3evUGWoVSJ9gX9
m/lcNuNbJOC9y7uh7NTCE1WxEdWIx8a5sUzO4R3sfa86/NiCUYdjyBqYIpjuJhUV
/He5crOPAzsnxjHInfTSzzJEjJQmIN3Y4MdBSw+XJHKtYhn3pXekbUN4n0uQV9A0
7VI6W7XrP+p8ytAuAaU+JgRZo9SJO/eKJH48yEg1qyrbgAW9hn8slIN+QtBXvsle
MFRHRYC8NEAXcZ2TRgFTDsLSrJRQeCSybu352NUFTvWvFwV/EhRD9ssxHjGwEH0H
WXJtOobKjth/c0ZBne46fjxStjJ2Yeg7pYb6v3xkBuo2fLlEwYBqcruYzsNeZLWc
HNZhSqWH9M1sEqY3+Lch7sMp6T3IyWKCKI01muBtyk/YjsiQY2i0nkM/bkuv4I0y
Ah7+D/WIpD+gNRiVTYS79YRAy8pl2ibes/jIL4I/tfve8eRQkQo03fWKufpFzzbI
4pGD245NLsQOtN2CmpAG1VV+nS+c9W1SUaGYSVhoavrxAAKxrgsSfDIt6HkBWa2V
+pLy5kc4chN6t6xAfbRE/DYCvhmjahmufr3HWtbVKjhiLSLtItncSPVBCzAW/4J9
m1rvTkH3onAxzoKzSyQiIlF/Z/0c1LcxKIrMPQaV42UCxp2fqEL7aezJVNT4DeWv
f2zo07qV7g+XUOUdzqD5XYDWnxsHaDAqSW1cEelVj55KYNjmlA/8291JfRn7YgDB
OkCJ5Vog6DG2s4OfqblxJc2cabTbQA9x0AxPEhGbcDtkEG4MCdlnG8s0P5ioK9kJ
u/2DZfRSscAXKthbgYGxLbVql4wlY9JblQgGfiWUSc7Xp5EgxODAlxAVaZUMMCdN
o9ZVtRO3AOjorYwnmJEqS+ap9IJqwbc66CGCjKMdxtxJ9Os3VQYTOjR2FSqjjQ7V
xhAX5IEKoLuCtQ3N9aHeW/HfsHMbT0xagqM5J+kU9LGXEZzPgdhVJbNq9wXl6keZ
ooYq2qqba4UZ0WkyZF4VB+ejIaxaHNs22J5rlG3kI36hcIUTxu3kraRYfDF2Co4i
fy53L6XjH0nE8q4lm1n0gLIU7/jiwpZn2fvWIqWGqB2JXAFXbYZ+TApc6esis75m
AXbgDt05wZMf0KsNO4wCLwtwGK22rQip1j7Nl1Kz730OQyRF7uoWkI9Ccn9B02mw
SNB/LbSjImbRJv42JX/cDYpfQq16XBV8bJcmgnwlfl4X7sTY2OspsiAdDKydsomw
7Et1CMTQV7+oIsywhiVqdDlRYbPZG6pbI6Em2I3GwPtWzXHYiDrU3sgXhdn7f3gX
aFWWJJQgKyDaB2gCI9sMJR/xwPXNptfqhP1BM4JY+qpXr4UfbIjs/6okftm2JO8U
R0kjCzgOsp7yJP6pWL5kh0IIVqcPjlwn+8HQF/B0Jxx11u9KuMGbavVdqxHgP6Wi
rxY6XA3Bvmacy4Go8tQz6ZT33bKvz2KI2aFJW8sgcvK4KQIDDZoyA65q8zRMkDU4
bvJnxHmnqN3YGFTAD/PuZZMfwnIqvamoJwD77blFnecfxXLcw3+DyuZESOLl7wvI
REhrnkfa+f/6l1MhO0j1qJ8YD+PkLp1KX6uHSBFjT1B1wR7zws/Gp1LyrDUKKvlO
/BEYuxAT8NYwApO/8Hi4Se2N76F9edAtb70t2Bhr5bWVhBkPjnmDQpO2N8h6un2C
DL7z4rqqKjpsRMGJLRVcKwBYXBd7xZt2s9eqByb8zHScLZ+/YMMD85qJDxSSBtTA
Kb+o08hNiRxMeM8DA/pO8O52tsQLuMJJHHRzlPllRLnjd+nCrcVSLd5N17i1cO98
GDjFpblyBuG4GmKquR3cjOrWNY8Eq0bMV3yT2dmQT52wl1AH/oYBgjoEc1TSE5S8
JnwewtTEHDXLq8OTtB9vbrCQ6KYluiY6NvAdqYNZuqf8U8rnD/T1VBIv6Pxrqd4h
0nPWZ7byrFWE8FVtOxay1nPtKGHn+2HxIekqwD1XSyn5DR9KaaDO9eP6z5G0Lo7I
cdbGX290Ni3Nh4KeTsnjIrAkpm7a5AKQgnxw5/tkSNOMK79fNEv7ahkVeORUHjWu
/E685aidvRFDiK02IJGsiex2+xrEFNDM1hBTyy82qrgKcBS7NZPjGghdlCewnxSq
7TtabnGspsqcErAddE8w1cfXV4TTgfo5avwAFXK4SjnO+dF6O1EoFEhpHpfyC+Tl
qJ04+haPX2bPxW1fW7SKV8eybglUU/IHEjtrnjjVOgMCZWvxciD8+73r+gw4qX4b
plDdy4Gg2vA8mrkAA2Vhvf8rYqExTyj7cDPqbTpOCb4pzVoa3H4bKw4hW0W9oVAM
baHt5on7PDsiZEdlJLa80cVOtpteYZq/hMgrRy3VD9RMs1EZfuC4UNYjWwiq6r1e
+L3L1JrrBUPjS8CEfV/3xMF5cf8jE1kZEDd2KMvkCKu4SBIlhu4ikSpKIKmGK4Rl
7z8DqDvIFSDC9UpcGak8nRG5kSC8uHERD+bk1nnnoFLolkIpDPPKbZxF/OgX5Nnj
U5KXvQrVJiOsonhLH1eZKXEfmQiWXnnANfBPVeMGPtSee3jlruULpg32xHFS2Vze
wE02+JBf3r4R21QWFBZH8zuZH0aX/61EHtuMJ2TFfQOxxASWpMvkb1ej6WOxO4zy
jvQwvrL4LkHx2vMY70FjgiY35/2F7uUuj1WRda0rQWfJfiQc0VIvpAPQOvSt3UzI
H1XyIkVD6+aBYFr0jYFgqf30/wrgPvYw3EHsyIiwDth9TWij1Jp99iNbrycdRt+Y
0tICrOETLSXKD+bHnZAOXE0cGc2XJdU2FBcgqwEX2Vn2myS1k8EPt8qq573rDaCu
8tNasgM08hiV1phLRifmhkgUBGicEdm3+Vof4Fsx9MafOMDTZpKP2B02CUPUtA7T
Uo/69sA4yN5+X2Em0cmjie3b/9s+uh8qADYPcdNITmo2iEnsbuEGm8N0A+20zCu4
oUSC2fGwFkQ5D+KnGtYLuBQ8Txjs/F/upJMwDdy/mAqsIsoBMEbVyvFHjTWb1jDx
J/Bs6zAk1d8E4Yc3vphH8sJ+WFVMGzbjjVBWjWuTkC7ee4KdHMJuPTunVvnL0l93
TnJXj9jbpZSMYpnnFNB538ft3zxlnmZMtpeqQI5xUUp6ouY0E6rJNhY/cUhQBSIc
mMWl2JVRLw2OQt6qC6rFK278p+qwBtE0rCwI/Na5pLeXoS0Sv67uhM1pgfme0Okn
BzqRdFurzNkXd3KXLKQpGQupPmpejVmNAySa0OYiJSGEri1DpeauVQrmI+EY0IAd
CYEsI1fZakwRlEC1B/j7GD69/OvFXkw+6R6hhviZ/hpOI7ibbUD0NbnmPG/36GHQ
AKKE1qxnt5qDEu22gWJcaGg9Xsi0srghZUYih8lttQw8Yq+gaO44q0loa0I0N4ed
SDlbSbmhlQU45qRw168uYgMlHX/CEj1d9tHMv6cx71dE/Qndhbps2Bw1O8NByH4P
3Y+N5l72/pQj1rhdr43dZ5ePEZV4xUTXTaExAN7VqePS9gUg2dU3jP9Ha8doytwj
817s8zBzjG92yzGRv3nfShnP2hmoRQe4t6KS2PlJnTpNZIciWi2BOtiNzv2qkeMZ
rnY2w/1GePwfbnOodQASiQvq87vtjtMrxxSD69a13inOk4B6cnotODcVin8r93Jm
C7DCxiqQpWwKi4yJHk09z0GosgoN6LqqlA4bjLGhWt3x4R4lGLUtBTHG+UtkBzAc
qQjU2sqa035bwgUEO4Gkk6yQiOUK6Oqdii/zqqiyddKtYYgT6xasdmHpOWrJp845
hkkbreUBJDrq/S2gfl1+F8Wk2FXJ5dPohxF+rOrS9aIKU64ncRqD8bzdaWTbaNY4
Jl7c57dXj2ZOs79rpbR7lP7UhXX2xO+ozOqfU/kn7RTTlaYwHvyXS1vgDWVV98Z+
wmge6kG6FV83scHPvcgfjK+F8MuY1SxHSoZUyCrostXMnU1uYu0qdUCzLqM8Rx5E
bOwcIDED5c+bIJN6ut4sd7qecVgTTfwsRvM2Ve+U8gnlJBVvLpW/3JKilFeVjoCd
pnpZOjNca3Z7P5Y936e/YbcYoxEtPyowTy2rFk3x7zs2FN7Anamf6ng90q+83qSI
RNDzb5EFvtIU6DcgYJGhXQvzktpkQLZEshA3ivRM/z6aYmPZzPEDylefJni2c9Lh
46Apq1grV2LC1YEi0wbUGVj4T4Kn0AI9+6tGn2WTev1kQo/5qaahkfoRTwlvh4lP
VDR2FS3TJBMOCCws3S6hqkNdTo1rzeER7tioGXmNSHFB2XnlOa3mVBePxKuHDXju
xzRdzeWsmmdj/yryqae8PTDYjYPNXIGDc2+YdwRxoPYom/2oJUTQB2iPkGRuEy2m
RvutMQ4CHIePjiooOUySadSQ9ZrEUhaZZ9VjmqGqvuXR+JUP4yX8h3wX5K5pjEOi
ZsUpCFyk4uOAuciZbyi7ws8TS/VfLe98X8qTLt2cxZ7IXpJ4jtragolwCcdFcVm2
TWT0oFA2Goz8yB4eJ86B3bO0UYjDpPIpAP0KU9WekVMoHZYDDhnO7S5ouG5CMHNV
IoQfFE39SK1GHSnBfvrD7nqp7fcdu7Q8gVy8A3bLEun0gWxNw05zKVOQs5KtytPJ
18ffhWTyWD1vI3KgQBIDo8TArDpfUOz1raMutMv3TmJ+6XqMyXDF6muZw7t6hGTQ
vE/a5UhbGaHR2qh+H5WJISyqckpE+Gx8Rx9BQQOnsiipNgsF1V8oVZ2FJRM+Q7ri
BZdIDF0/Jk4XT3KfA3uRBidK4HKVEbXhsEkubgUtYnCokJZmLGfrBM5s/DALUelH
D1AWpHfjRd5ulf1Ci5QHPS4TeHYPJQBQzNqve2LV3IvT0EjPz1d5moJG1f7lsfdj
UW/YEAy2vE823moZsqmzmUMnMmUe4rKrIxisYUFJidW7zAS4sHmsbilNzZCmVUw+
dUxOiHy65iDgOi7mR2Rgk3dL9MCFDvCZqISH1D9UFsxDbp1W0yLMR8YQWAEg6Q7r
pftMx3LeoNwYiGasxkPJY3FilbU+9eOBrHiH7Zt/OLuL6sNLmD9nEV2fqH/OggTt
ZnQBTnnB9sgztL3yu19X7xm+nHzfLyhO9NGQaufATLMelueKTsJaLTgyXZAKI62C
RXcpz7evbgeAYeNqs4+9T5m6aaUxdBxXZuzNLizyvOn5Uap211VnnfIctq2XAgS+
UTztgoSS/rV9s2r5z6purh8dkJi7FS7gQdRl/kw3JGbDOpeMWbtAq/7p4hF85Vzl
EiTmdrNH1c+sbZcLH5n92VgaThxV/I73rjv1AXVgTkmzN7xOZa75sJja2AGc5HrL
2bwwyWy9Rfj6NwzOYg/E4XBS1JtLii7wGufj3fYsf7YnPXlgURX89P7n6wbHZ2pV
iMyqJq2ynmB8OxeE1FJk7M4lVu/YrJOH/YQ5BWNmLl3LhBRFFOaRWD5uXsPwilDR
5UJj+0mZ58rKseCNbR7vj7TityZ60vGsRppHatsrnEtV0j4yaCjYigr0ZKZ90A6p
F7xuRvsSAgnqx8fS9lK91EZgfcqkPvVzH58qii+e9MxuICS2zgmf8XwGDZxMUPlF
oox0Q0SDyxJaU7iwlsqe46o1t+/ZsXYQoASaGN4gmJfKUeN7yxCMEPlndpbfM+F7
DllfzPkT3n2zhsVMAC6/v8Q025tMBRHzY7H6jGiZbBhCJ+dWBEC8IG6e4EzLBl/3
91AwZmksiT19Bw4qGXcfgd6F3xT2kA5pUt3J0wDKMGqMmwpPZ+jguBMWdW76/ARt
XrFUGtVmZ+lY8oKfgRz1PxwvPJhrJwFcdhRKLhGyMpePSKvB7zs8PMcLjWKW0osJ
I26jiS16I7NvnVAElrC1RMlo1VTlmQ2d020hZYdkQgK0BCymfoESiu8n7FzP6nAg
Rcc4CSpZpH4cobfLZrD5Qy7KTp5hko84Qe2+rTTwUB/iqSxfMmW4awX0YIKE6UuG
Nt4rAQIgB8bJY6G15UdgiUz6+gKwW7VlhaP0HimZysYRwP820N03QtGQDEZxV3iK
ZZMIbCdMfVcpJFIAQNPnU8WZCNLh+r+Sk59MK+PSJGnbdagiBcDEtYcJjCDERu1e
qYo+3fOyVwQvnv9o76YGhnIUE5noCu4UYwAIqaKC6NoiyJ55X18VvZURrFOkaPHV
G7M0nLcLCXNcJw0toUBM5CmjA5/KZFYr2uuQRGe9YIzjdnKhh7OsXKE8JlVnNiW5
wRlV+eh1GjXAt4MxlJJ8STYNZK25C65RyLjUe6vtG8GVQ6tuEFdmm+qSf/0Cl9oq
/2iyv97YxolElJ/v+np4Zv32buAwIgwshPpeshYlwPrzcTNfErq/g1qKMI/HUKqT
lvm9XKMNykC8sJSSXJ/M49Qs+lkABfs2VqY3chUXF2H4R2GqsWC6t01yWEHICkz+
RSEmMxqqN0xlg+LYG3GxtFAfWPL06HAup12L8FsQ1l8spo8f7wO75cDrod9V4y2l
SUyzXsrRnBA2UC8AlpaAQ0P8AfpSc4Ef3WpxAZB9togb5mGoxukC8GukfxCqcNP+
LnXIv6UO6462Ah41IN4TYQ2BWdvY5zMp6fezPXEjWCvXolDytTk/FUpR+khd8ABn
CIV4UTGcTiOJZr+r5UHpE9hJ39BsqUwsAZOzcde/XjFKIvcN4CF6g19+p4EuJIs7
P5nTvz+DGmayKi5JyIgGAWJ/S3kWyDKJqOvZGv0y5OqWAys+IAmqXOHEi8HchZ60
Cxk2dnnjRbwEVrSw1dSpy8hTM9jxlo3/F2D6g88FBwef7MmWAaPVFG5124wJB0K4
SSNc+Dv288p1V08V1Eiv/tc4dRjs02eXJllP4Q/74QhsczCXz5/ODZT8qpu6oj/i
Bk+Gmky8KagetYgXuQJuiXPzKPoFKlf9YOPjOuyBQcJgChgsBCN+Y3ODxgaIvyfv
oNyV98KfvhBrCeTIgETvJAngZmU9MDGA5q8dL7qDrLXf28iE1w7QHe3gLRD0TMNV
Psk9bfN7i08539JnX6olqGDViv1AVQfMEDkUZL/tCv+8XWe7CwcwMqFPnHPJLOeH
OUuyyu8iSwLfwtvMeQWl5Lso1ZrMnty++0glnXK/9zOTmWPHTkFjIFJ4Bl3bz0xH
4tScaA8n0ebkDZ5JRQ1oRfxmU0gIPk3ShCGwacjThLq1L9n9P6jCHLHtBlTbqtM3
gIXSzT1287aunqlRzliu+6aAuq1Rmo4JTb/0AwGmdCsfs3kc+UzpTOkVMnXoEn9L
xa8vGaXzwLPY/32dpd3/t6IEHXLaNqYB577X6gpORoweBEsVsNqG8wvfDzk5T+i0
eOxT+R6KGRECPmI/Caf2rV5WJ0S4x6sNwbx4qmq61nthcm8SYQaC4oA46zUmoZ9F
/sHIJLBF8unhZvYGBeWpPWsKWacqUCbeb106zgGPTAE2GfvSMJIBFFhMvfYL46KB
X9MsKi+hsMUryhhV85T2aUlDOgNyPDFg8t0ooPdbGO+ZqiDom1L5vx7zQEBNi4Xn
qtCloJ+iJxD1ysF2bav/A6hhWM1J+E/As3ld4iGfnk+JVOsUukpHFCVG6efe7xil
qEuLAyuccCOdYjCS0Jj0dAKOPtwnjn746j2P16cqmF4yRB+9H2rNexXxvBNH2jAV
Z4GiqUdUscywpchybQa2XW7rYnXEKfcK7cN1GPZV1/cbmyFcGTvGhW0SeW7Sfvtr
fz4ueVQE3lENp82vbFXvnm1pDJ3xZ8wNFCcC8bnjyG8L/r0caBxouOEpJdkq3qBX
wyLY03rwAdcQH0Kz1OSTqVrF5lgQ4fG02qgqJ9revg9wXlMYhK/6iQAzLkZkpYK5
XiNQJa4mh0CEvilNN0bHqIlLW/SnkgFsgNgk7PiylxdBYSBPy3t1D9E+AeF+SWK9
Vy4l7iDaSS5NGF7Ohqhstq5ccnYgVair65zH4IlB6vebxIO+mJz0G1Q5eRkgo6bK
aZMJ0YaWRtcC2+kisjR92vaJj1ccZtgpIjmTHHJJ0fy9xU+jw7lMI0QXpdcXwPQg
13rGCQUOLBcfg2F4noQ0NjqWIw67RqO/mrQQAmx84k5WFlb4CpRgEwaf3zpUEXgR
T+Fp9JCxhk1P+FA0RZNvs6cSqApCG/CBOzKlyYDO/hlNDtC8fG4/RDHJPSrL61DS
ZXJMHks75T4JaR028BFVKK7AX06A/UNWPyGy2nkyCbsWFoDefCa8YaBVv3WDD2yr
4Zs5yJRp3lfObev/MC418nG+EqEb+Tbmvs0kBn57RwRPPgid6ITOP5srZj/jDsi1
2QPyxV4bm5koFWkjEQrlMYulRmyqS0zhoybWlpKhToL4GwQvu6xKbqM2lAV+J1A2
Y1biUFVkB9wVFxE1Ai3P7kGrkbQyne5lVzpFTaZtlij34kt4D1ElF16MUVha9LWo
YNEqyUz9cr9ffgjF/GAmX2nttOkcdi/xzJP/XuB7HN8EEf9UIlMGo9wAEdMw5rDy
+hkK8KqcBaxBjCMD8MfxJKDg+OImG2SJy8/RuoXOZCcT3vBpFp2ipNjflegk0v4d
+rSJO25NkfdoduxYcO58MiVRsCFd3TD3qpQmczrjYI00Zj9LURlVmckTPTrY77JW
z/gQv/b1OKrNA7BAxDzsHV8tUJ2V7C7haYLAsa/2WpHR+53SrIS2QD7catZ1fIwh
mLuZBmQUgXGuah0NgKQVZGrlooAZ9+xqv25q+F5Hf2atzus1F1p5QMxF5HaD83WQ
KsSBrTmvgl9TpQlknfqzDtCjBY8u7jrNvw+iS5QAYW28H6nRwf8mzb/nw9VV5O8Z
ZQcurtCC2gYeOWO3RDtt/SRKxitbPV4nqQhSYHN4vlRhTZ7VAl1ZbhkD2HvWCtIU
FKnhxZo30dtlIlqzeBuIZg5UF6WJoDrC0CdjXAvZWV/82dy8Ib2K4NBIToJhgaoH
poL0LcDV8hDzT4uT8fs7vRmHeDMVYrBhfXfRMcrRq88UiR5MOhyBG190bwwu2Jkq
j7N9neUmSmxK2uD4wZNiXp6siU3cjuLFUP1R5m/ljFrJyiSUIXOVrO7b+2jyEJKu
iPgOdJ79ocNEle6TamEUpFG6nH7EfGfh8C+wNa/MN70TT/SCDliAWN8pJDFm9EP9
rhiOJnJ61qraoMmigucHD4OHGGYlH6r6RfNX+zNRRbEl3l/ImbaDkyC9n4EE//yC
DJHTKDL45XutIszUfpGCnWr4XxbAZeKm2dvmDPht3XyO6wGIN62aOgNNyel2L8EG
p7VG4/pdQN5I7Ptd2P49TNZLs8v/+lSRGkreiv5JxzUAdgIURjaegWYfxloXAYEG
YhZ9vilHKWnhqd43XaO0F0DRL1l3XofPNPllFBgvaNOPG0YMJqxfenCypGft83xd
7kS9qMQ6SVrVVgt92t5LXjlBnQL0GGa7TuxFoGq3d8L3VitOW++B//GRM2YA4NJo
sf9GIil5oO4Sl5fZmj66keRRtNv/PKGup80r1aluXuP6hUrcnpFIEjfPOXTuX2pl
dXz7UxvEJ7ExD90CMQaPy5mTLL5QceFLAbWKrvD+mlT7M04EHQ8qfSWHo/vSV/Tp
WOqT8yLNdxmzbm6jbmopSvk7I7IdAfqnuSYyjhouNA+J6GdaeNfM0JJ2eTOk/sBb
XQf8NROOAFpQW/ivbWYBw9IAg3U8aUjpW9PmGUyb9sQlzrMSpuwEnKXkgmNH5bII
RNzAxem9Pez/S8a2cBdhgEBRs/FWkbPyind2D8S6VMKTTY88WuCHXiVUnbBzPd/t
erpnWukplhjnZXlyXHpzAWlbwf/+t3+HJieUoPwGAu027O3AB50alrnwo5CFRYiP
s/na6r0DSNDS/QHzreKI/GPCg/LtClagrAWFzv+y6sSia50CXXqVkwP5dUQq0cNK
ot4RX+Rpoc9ZjGOEnl8pL38EHml/MsyGC5ILGqz1IBCzpskj2svroUVAs1yIvmol
NUe6GquoVwdaDKaLV7s8j2KNUyYUfmUPaVIaa6VRxfSPuTTKKEDiq0Q5ws3n0mB8
Xub7Fdb8W9DsvVLeA8T4k5WD5cGV16jhH0p5c7mtTmw0bG3AvupPuYd6aM4R65Ff
2D/pU67ZPNF3FdHYVFcsLIrEL4D4yhZNMWofB1GFfW+s4B5twZV4UJGRl9E9nJ5B
Tm8yGjAV6DP1nHpEZwQKgTWAm7hlJx0BIzmVuHKKH7NULTziEuhiVYY+uOd/VBEo
QfZVEc4sDkXvHPGKKlxssf4FJ6fkKzm3DO+nbzamrsemexEW4j5nOyE69xJOL43S
tJYy3jMwZT5FvKy+25kNkBsgZlQffGiU/ahD8QPrJJ8M5lVtO7MNAvraESnSEG6Z
k/UEZhheKdfdB3aF/UU85IIZnPG/nEg7UcyaTLiuEfFNkmtvkmGqFsP130xZ/7Ec
8Kvy4rssbvGQFYGQh6E7eg9VRHSthcZ7e7pyKP9sHH6/G/ogeWolwt5Sbf37cZXr
kIUFDcUGRR42iDv2yUJkAGmt9RPaFRdcCWl20BQNqORuw1FZv3MTsU62aN1IoGAs
Wr2Pbama2bMyVl4VR27H5PWXS4Od/kkT0UPmyb40eGdxWr2MqfVje49oQki4b15U
6/gV9ZyBQqZ7mved7r0c0ahmz/sEdzeC9EfR86xccOcvNDERLJ7LwUK5NY1Xxv18
gCzaOIfW23lJ/q7LtkFiqgnkhHUzA68IhWT2ppb4JFiwhlChGNtulSNNlUo/IqXG
Ogfn9Ypw0BDI/ApgPwFew0zSBHwvzqOBZNRdb7krKFj4VR9xg9l+YxaMLm+DuKLP
dvbRHvw4ZpCl/yqimJjfDA1eezTDqq8YdPT8x6uKRKe3k57HwqPFwk6hyaAlAhmk
MuA5wVRPOVoSwZThsmSuUKfiUZvo0iVY+OKp37MahMEEtjasZh0ibNBkywtRPbFT
UHNWKI0fboENzbilUdLCgOyXv1e29DYn5df6N3xujxsgtY851P5Czjpv4v52yBF9
sIf78b6X/07cEVmg2NC2m4z4hLHDcHZyea83vg4S3pdAkz+QRKrRmFGiOD1QSBcP
UImJmkscD/SgfeJb947RV5GlC/3OjnfirUkM1HcfikVjTuaJoWj3pdoGR2u+Gdtw
ysJvO1ebkvflZdGnBH/t2FIYq8UkqWT1T4pQrT8CxFhSfCoKkiR6iSzoZoa2l33Q
37Jlo/AqnmiGyzXjTGgPtIg+uZvsyprNJ1i21hEfmAt9OotRm0VInJSDr22ADgQp
9FcHGu3yxl8kTzWKd+GAoeuAukpB1HlOmHRC+FhlKfErh2nGiX4qZWOfj6crrhjQ
ACg8H+zh1KEtXneQzZAXAakuEYEgK8i3bV4HcJWOBZS0V/z4JlduF9+hiuXk+xVX
Nl6BwQpbkmUmWLYRBVqahAr4pjbhC1tNNC6qfoMmqmJS7qu2i0V9iDbuI9TN4U24
y3IryuP3hRb8SEh6oXFYM0fEMPoBz1WU3DaWvCFc8OQXOPP49KEztzKNnf17HLDO
RdRB+92E/EqD+oO7LvAaMSjUQS8qM2o+vkGtE2Mva51jA8m6qlSdrNswW/DgkjDf
bfQM/2Z5C7J2knJUFwwEAILC3Mr3+vxJVOCg1cPZgiR3LLZ9VxHoPydu1HENpo1k
u+ZhWjd/3SICsHuPv/dLytY5BSJYWG7p7UierV39B9sWVA2P2Bi4oTXW1X0VJNuf
eBDnosd5ALttIRItT074pJppOhuJlmBxWj7DNaY3FAs9lb1KntPheHLy+6R/mNyh
lpzXQ0DXCLy9QtrOglL1TxzcNPckL0jpQaU9fxnC/vHOqBuLeljid/S2v9n2oHCR
5gfnFPAayi1y+ZeQSt5t/hnMqdX62DfmHAlO/0W4VtiKb57/VXX+NLW8d5uAC7MI
2d1RrK50TrYf9BSD8jY8eyTbKaBwHnya3UDoUmaNQxuskfaa6O3V0oasOfqvRg1E
GWGjvKsHJm8n85AySTGAG186WshAswZrzLY6B5oPxk9PEEzfufMYVfYQvgwL0S21
BUP6MYU1CVJr4mR8cMnPs31ja7QdgGPKeKDqARrRzmz5ZSR3eLzguweUGcQiLxxa
oaPJ4Sbw8cVTKK9RE+hkBuJxa3eoDe0reaNiFnXsX2TocR0JliNbpnKCKcjts162
hnhF8I6mJOq5a/0I/OMix4jQjewHoUGzWrlKXaJUFYEZDmQ1019Ea+Upy8VWGhRL
hBzom1rYstJ+QX8LyGaFIkBoqopneevjgsbUEpnQzVNeH5zfN7sgKJE0grsWntsc
xP7M3YK0cKHJetD0CsL8Y+uFxFrhqM22d2q0psj15U5r5aMFXO2k6OVB622owtzh
cE2pc50YWYSJJo33syWatQ5hyoJ6MJa+B802CDpAiEPRckf7GvR1mWQMf5Tma54x
sDofdA0kqv8oIJLvRqclYbH4fOPzbhA+eHuuLM+7iHqd45oZm7iU1JgkFs67Kp1o
fLBJaa7gbslgnhfhB42IZkVWsCsgHgNn6KsncuU49dEctL9fIOZ3C1qGiLfQnvl5
W/UWU1x+BJLuHdlln9B7ELG5ZpkHnZfRRnh5yS1gDYGj9HJ2FNGGDZkd96M6J6QL
e7xZh9M8XSN1TqgE2YCnevxCfbw2t5ivPsgq6mnf/4WWZN+/jHZBdFWlMqUY7Fe4
MFynIYPlU5m4ocl1lJe47o3WybKgCdX5Bqr4YY4Y14/DjZufYCwqUSUnFH+xlYBr
YSkBA6XIzJe7rvpu2lziwEPqX/n6ji8eL6Cm9mywiKgmUrh/GRPYObINpDT1A9Db
C6pvp789xXS3b4SzpLUeRrB5rw8/MumhSjuyrbz95PQcDk51BQeK6gbnOhWedG9q
m9RmTPkpPDdk142BCCQnOrB8oqgG1AvTq3nBAXt4/bOsoZjnQ3663FnT1yD4eIjG
87kOFm6nPNuH3n8hJeqDnUqQI/OFAVcrOhjAVtAiB1HI5hAp8ZwjTtWzWpJU8Qhf
lWvO3f2hA4BKdZkinS1MtgIHFWrZRtpBQmj6ySzP1AtOfXtb7++OAD6VsDbuLfCy
yoySsL78Ozb029a4xQrnkPDzV3UdAqn3yp1rhaqcticLOedNOv94jXCuRhZloNMW
jMG7ld/9pc8XelSs5IWJFnZ69og/Q8DO3QN922VwwkV0bsNm6NpLIQ2WTfyKRXVq
1qvoUri8AXMXyEGSLvpNtKQuwUlNKmuy565HIZJPsRupCRIFFMsbnibQ41S8YJ9n
VS3RGsn8P26a7S5tP25xrp3PhC41kDDVMBxB1oKxUnh4cKvjFZk8v3WLywzZSSpV
n3L735Z3yc2F78Uy+vlY6QdxkTiF1xB5zXUKUaFWtxFbIq3S05qnRrY9B9BS0hVj
aIRJ4bnJ4f1YrtA9mYG+aGNtEhcDhv8HEM5wiRXYyBoMpeT1So2V4ux+l2rgxt4N
152G0QOKO8ukR2bp/ZRI78V/LI5Y7SD3r/GcfmGcp0aygudg5O+0JzxcJt6y+u5L
ouceXPD1jZG+55578NiHcp0pf8Lp9kTP2MaUApMg2O06B1+BZdTbbjYWN5xiLqrQ
yjgeBZjXG8Jt9vSH/6TvzEPljy0w8MsWsjglgmGDr/wWud8Ie0bkwbgkI8uVIcw3
bW1JhO87++xJDV3PGN2cOnvgm5iWTbWAMfua1ECqK2Nja7cA9Rm1Bj+0biqythnt
AfQHhCkBSH4yAI9lQfXK3V5gs33wa8+oZrammJWhmCOrsrTBPV0ks66ERYQ+JGU0
RGCRbMQ6CkP/if9zDyLwJZTzPKFLlRH0k6v9NNBVRbCROVA82OW25408/mvK/8vY
xtVt8RTueg1XVRP54Sdu/mfLx3uErwq6er2otyYihqIUVoxQkZyEmDJJK37UkNXd
8oAOa7LCsUFroc4JGEp0uHCbFlwWV7bwuI5/a3uHmk2hTcPA67vck6m5nwHPsv3H
XknEnM8LmlXgIrzSTK241PCtWKy7LH/bSX25Mw6xVbStzHBUhLEU9iGpDWobwMGg
QLkdiOE4qNfGG/KLceR3+EtTuTlctwptRMSIpwI39XGwzDoE0RZ2WIyD2VD4bjoO
1tVbo8ugS6WeIWbFyTHIN3Tzw+pEupGKJVsfSO8wpBeRI22viyCaDu8cRczFQzpR
2U2m+7Eb3fPZRhirjc9KBhcz3oPBcxq7dGK61ILuZYUcC14YJ79FO2n7dZL/MCmD
HN5pJxAYG8a741P5WWLCMLf0ZAZEGQAIk2hg5UHNPvUbhtEc7WBygdKMrzaUp3JB
wZrTAvUIzRuCLzqMnlzw8xDbd/xieUIQh6+SlEY0iCDTKFtlVmZfmXnAWLRdWXad
3ZQk0qH1RaCmPAhGkWHrpHnxk6jKwEZmLp+EOX5534BBid6Sz/b1WcQ/wt4FyrT2
2qUkuwwLwdOSNO4Wuq9+Fn1PX5dReQA9NoaDRpruSmcpfNtou1LTawuOAuL2CgBd
XsDNLPZMQko3cf7G8FWLYhfXOFBrkHdsJ8c6iPlJdgztZovyItGb4qZXmRuzwphJ
4CV2EuVVTkIJCQAD+L0QD+lHcSnBPjbnVU9XJLiDvcauYj3NohD6GdG5Zx5tZvar
cQ3hD9xEHeEYjFD8C5X9QjFnf6ynkO5lGlsULgS9wUH/X3aQP1YilIC3zX+84TDZ
48kRWO+nqsPlprW5HHpqjJH2xuijcdKkYFjrpCR1fN8BTd/EBDSOjvmJRhrfk/Wx
Hu2nIqi719N9eTtTJKSlLZI2qmh3qyqO5q3zGP49TlzR4GQONL/0JHTIlLDNeKFX
WHkg7iJU/AqAZSwBu8TQHD5EkeNwFRROJKjwX/1tkTPjqGwXhtMTfKUQIGIMhe+1
MYrEyklEh0FoMtOQyUfLQMZacCuY1U/y8yNAIPSGot3+M82TN+7kxXKamGOYKLCU
49jYNvfs6+HO1utqtTyI00mNLDdqU/+ADGvcJaPFv48ha+YIRd1rINj+siuCtOd3
NG38G1H+c/B2DdlxqEVEZBseBS4XUrO9Cc7IC27e6AnaCDJSznvCxcdXOGo0Yyjl
A1cKM5iOCb9RKPExpjyeTy4NsADcTWY4HNww5tdG4e5dpNSzhUpWqDNUZ1tM4uSI
NCShtdraaEZ4lDB1Cp2MgtDTrgTt9z+qwgECIVUrr6ljRXW/i5jrLoCJqnK8DrfS
kymoZYq6Fknb/Pb/eBbEY2khZgMekjUBSOO4JIQC1ZOljB9WGyLAVLY9tP/pDxBm
p0JBcyHdYvgaHZgolUeHUbN71yF9+OvRhgXv4I0ftSr9s1Fb7nLF38L12dfnWWba
fgdKyf0oranHWxnQa1aqCOzK23kcJNKeyM9BGsYK7R6KQWuj9o5e7EFUObBb+a0E
5HKTTuMo4ic1qs1rxS1/9A7+JSz+9uAXUHWC04eS6aOKVd9Gl86gv2hPbLI3Hb1P
9nrhZ2UDgCdN82UxoTYAIkBJDO5bXiTqYwyhbd5Sm+r0RlfeubGlf3G6eAJQcusM
Q8Xb409RGUeukXSWMlfX9tu5iIEYmN7raRq/GY5LDEruxRQ26To2MQ8mu//mC14R
He6uzjTCT+BsgN2p4u0VylwYo+N5KYm0Yl/qc2EfwTkTxZp59V6ILwkMOb07TLNk
psJl/vlZ3ve9Ig36yRHwZazMmRJEYc7F1CDdbPOUgaDEdP7wjnGhMO01pg4rXTis
63R6YpdjHxphj4VN5SSlr0AQhHDXwx/upkfyEXvjnw6wyJVwxL1mGknTOngn2rEb
ZTcglIb1kJMD1SgpqNYK9UvFERp/iAdiEt+4YPZUst+kSFbcXnk7iOBl5rAVPlZm
Smb8fgTn/wWDV4mGvXfc9+dVrdR+DMEy60SJtw8TQtZHdA0XSnSE32EC/S2ZtfJl
uU1s4wJUdmgTTEwrOhNRDwVuedWfQj2l+vNLNrexu8PlZ7CuX9Wt23R37cm4UGA2
Vj1nJXLyKJaFdJN/y24s0JXxTontImyIWN27aknqAaDjPCQTepvkxsZ0ltfLua7c
u9lp/KVtmSvw8V9ns7UfDusKVUrQpCan8rqbVLZ+/fFUWDyGQPLoZJReubkxpBLY
CCNtaWozuj2GrHmdz+3SO1nLOxaOtYsqzDOpPxrwB5g3dn6Nolr3G+3zwJ1uWgBf
eBmBKF7WMz1uYT7cNVRw3kliQNJ+SX4JTU6RkHgjkUIQrt/2BnAW5y0/g0463Sa6
d9/DKdsR0q0/Pe2lZM0OVm7sN36mWMLIJ6N3dh8zA73jNGSeSvAa/sqB0ON90jF6
76UoPK0Qj0RhkRUrMhwEXKcsXuuxCNnKyPJ8GRRBqQNT8Fz0jB1HQBmOEe2sSpPF
e+5u3SlzJw4jYAxHDnzMVJ12Bv2BcqX7Pryz3HQHvwTif/rV4zQnA/nPfH/EIVUQ
BskNfQ8prmiSwcJiYh5y2PMP/R++FsunwG8CEo8sgZTaoQU2rfOIaHXNOWfpEq0N
sI3n/CfgoZdSdbQRrziXS0qSUIpm+nob05TCPVonNnuZeyGbAtaAL8lftJusqVn0
a7YnqyzTi/ld8gtlJp6rffQgFhAnEVqtxAxVwHN7nCoaqvjo9ruZaauHHfztfMeb
7O+V7mzk1K68kfqXDQvp3DmudxcMErtCGiEHeWOsr4iI11wgemjpTtPe8GzENyaY
RCXJTN4oMXp+8dKw9V3Tsmsw6R2MYDf14Si/wf/D89uAZnROZloIHxbf/S2WBION
fa59g2gTdsspvwVRa4gPVKwTMODdHyMBVcrK7+IXozJAwvGiaADf3le7MdbVGFPj
9JFOw3XbchrWe0k3fulcvWn2QTkVut6WFbH8GP1iu26NsZc5U6hYt/qrVICOYw2i
A4OdEESMGD5sXu4KqX/TBvATNeEjGP3DnCpXqusLUJW72zBPS6sc1z2hj+egEoM9
3feE4JONycr9eFpKzQS2GKyyAacf5y89wykBeM4tmsgx7aHPWod3/Ps6wAuCIUTo
fhyBTJ8Cm+cQSZDHAtc7NsmB0G7NlUtyQ2q/ciewFHimzDkQQgbaeQHVP+KEtqZD
et/C5LLdODgDafIJnqCiS7KaJ09oKU7f0H8h3ho2PFQBOZoLVSU1tjOE1z7shEgv
4JNAMwG5WXFDcirkTdthYeCCR2/pXBrsdxcL56sLVJ3IafzAGrqIOs17PPD0/o8y
X3MmfnmP98iyQM5elPe7e7BxBLPf4Dvq6jSsbtJmD/WyzcMxYltsuGJziFT2VjJP
69vJguPw0mWLdWSKK8A1tdSUuLKDZZQy9LyLAWVsqJ8NIWg2QjgqQLTfA5wenTC9
HgwDEllzyN2Fx/ETajPAQSVTwnDR5gLyQL5AVBQX0FE2y+98KyBPgFyAZdwPm/JB
x1SndTsKgUTTs+AGyI3XX4bkttJk8ow2UVeyh8tVei31wzsW05sl3gphqT8YE5uR
pzRmtJ3Vt7v/EfwOBfNSrzp+3oZHa4ZsxndRwGd8oABSbEoZ3Zms3R7LvyW6uZ6L
h6+mzdpGyf9xMDR9sNryGAPCj36vDUUvFoyuYP4vti/IInfzWI2WhBC1heLq9R8R
rlAiDxZeJhpPZRuDId82sgmh0IKLC+zsPAOMKlk9Y7gffDsf41Lh1pVKyzbPi9vE
Ep55yg9FTFU80mR13xgwg1TuO+UHmMum7OWuvgzVCTcl2eWvh3KU8N46IosgVUVp
DWcdhyyvbpkuBgJd+7SSkjCvoKP+eFlPaEzWiI++LSNPWailZGqopygAy0MVgVkU
/9W2U+HtDV0Ij5DnhIdLxsfH/dhAC4EMCrpJxt5T5L55X9bAjcvXyIr6ZX6+jOb9
cJTmNp+0M19nan4mAr9MEnUZwBgV1R4xUYUtY8KRkDAFrK6chIl10pBSW2D5WKTw
0LqtNRt/nvtX+vIOxpa034Kox9ndYF50pR7uXrYrZbzlZcy7rqgah6ABB3JTJw3b
oYWLi53BOJY964SkifMGS50J+iCChV4eZXaT+OVtKhxB5Zat12n3QGB2qcrDFGkU
FtFN2ncHK/dWhPO+MmJwZM7QbvOPBFweIH1k+WNfGN3hwIv/Ldqps86/ZgwLR0pS
DMFdMQYd8X7csPgTxPhGzaHdm6jtY8r9KUSgPFK8kbB6vI0tG2Gx6oIX5uamGlXt
w13DIlySw7X0cER93KsPHEMLnh1JKfLhuBcSn5ZasacdG4wvu9GaxOZO4G+3Xttc
8r4Bv/UkJfrY833xt2Lf5hnVoaLvfiOZ3FwzvuVNgcrrTZogMhYU2bKmTvoxaSOM
ExG+4qnRQzV4hKJx+GaxQIYnuN6Vuw8HEFNQxtbmczakAeQ+Jweo5moh5WWbUxA+
/SURbEf8OupLm9zrrNUwP7mb0Zf/evMXpJHRztexLPxV9+fhr8jjzyUmhxehQGcZ
/J5ViNUCfnK6Oa646/kvC1MInBUdp1/68a2EB/2sW2PacBwmY6peqSz0gaYgOJYH
eGJC6KIvJiE22x3uuPzQEDPgtg5AL0QvgNnsDPrWybPZT1UAgeFkzjvgfMioe1Se
4RCRz9QiJQOM7ZW0WUja3Ydn9eOCmE559RHKUKftLyxvDrxgK97UzT7mDT3qZCRV
QUAsXmoyjWvV+VArJ9bOCzLNzGATT810GQRvM9fTpNndfnSL1JEUPoo8H87llBDA
+IE4+78Gi9tPHsjDRXKjtaocs95+yCUKkRTFB7SMcD2stEO3W8ZnEtNh5vX7piuQ
vCcN/AYZhGPMGAxA1dRa36qPmW/Zo0mm56oUzkMraYuMSm2QQq7bm40bLx0UR46r
TOuJxL6KrLARsD4YG994or42LFy/Mkd6B6KFIHQLSLD2tmd3hWDJfEXq9JGnMvTv
P8Zix7TiyS9i8arxBlFtEbZqBvX5+6hLoZ3AczJ+VvhlZYgeLhwffujhhYfUDBG3
8zX0+W9ZJxONRjU0RFPNJiKuRh4hBlBA1rheCfPm55EH909cJbe2RZoFTT8XLFgj
tqULyNLuHNKEDZmWEue/a4r+ZP1vv0pOPzTXYZIMjnLEc5TXlbLI1/yLrrYBWeYo
DOTiOcTItaNscXQH15KhXyTKAYWlTQx4TwUsUNQ9YWOZOzfBqEhI8kcEDNxEvwE0
pXb6F/LXnnhDzf3TZut3ZsnksJtme/SOKCNJb1BCfsT4BXxe69uW2d2H1QYJKh40
muFSpeEfDucnOCzct+I9Lf0ID9BaE+G7fapar3L8fCQvmXr96t5rU+0/crRnN6/i
DClgF0LiQkBh9/5QIt8jAO6F6UZZBX81pIZ/67i8835/JXugyzsxWDihI0+TLDRK
Jtgil3ORThuOb3qoxZgLUBaC7piVhDhFH94oxreMasDUt9yHy38v3mbr7b5JBcbd
Inj8/roT0YDoqNY8eXP83T5EhfxN0UfusZhDaZvb5zSe8M2gCTxOU+CgJY/tiTWj
kElyK0KtwyWddT3iXHY5aFPgOfPDshmRJQ+PcyouXypJtVg9m+bfPxF4BXYYjvEP
2MuIrcbCIufENo0CcSDa98pZwDtQeYSQJOa4sBuBb+NlAHJhmoX5lBuuYpD3RMyv
f4rhCEZmZu45TrItCkER+kPlIjOdz4fv+O0ED+Lk59qdSDg0v3TM6QiZjONgtR0C
f84pTi7iRlmCuE52TLHInJlXxHBdj1q29wOfkuOrP9g33wNvfcpgE8YECq5l25RU
oPkBEnM9LyGU1dIxPvFVvQZWU+8sBFnqd5nG9uRCUrPUPr0ybg7LcJecm6BFxz/W
lQvRA1G0pxrNxOd7THCCyiuQ8ZVtk79GBDi7Ncb4t/aYBuFWahC8o0euJvD75QGs
JFlCJvcTIMXWDLAuTkOrog437kchMdCjp7txOSzwJI/304ycPB7/Ylt2H7BnUEZq
DkKl8DUc8MypKabhTx32c/6gaYWQAGFxLf/LIFU8xob+aTAhCIabZrTMjGWRDshW
GJ6gDqe/ciSNUSBj6SKY953qz581rUW+ZJ/P5q/nw43BWklJAI3wG3+CdBTAzQQG
VfDOyTvZvez1469jwixex/qWtq/SJ0/44xiHYqXmpoZEcV5IVXnmJ8LGvtTmjBeB
t3JfWR9CzZRT9LeywnMWRCP0hA90lwYv2j+zFbRvZN2uQCCKboy5xL0dybssYvxO
rpSGZIfRej6CqnIbixljXOC3QWqwvfpJiXSAiuSCvn1amEXCWLzBvDYPg2cFnwUM
FsxPni1h/FB0IQZs6hhF3er0aOEO7o/Z3cQAXzrOsLfxwCtkQQPMQahQjgV1Mi+k
Cp8GIWZIWX9MzptWrJZLlKit6PeVPxJpjlzrdKC/ucA2dHV2GmAOVVOBkK9dWhDO
GwvpK2pwIVczT4GfiaSsi2GcZsjzm7srRdLJP0iQK+FtlaQvAE4SfrW+EljpsvF+
S4tH6y5KWowY7SpFO7XtqUnlTDl5xPqgQoWj5ygJOw+BXTDW4MOYYHyi+p2dAsTF
Yz/DmF0BMJrQR/8GgOxyV1HpqxBVPK9Rv0Vr9OozKr3fEHh5fNXNgD2Mt9AsyTav
RiZ4fkIvKYB5fQ04ddfdnrAWku62yVHzVMvYDM3peJ74lO4+BOWIlcJfhEzLC8ug
SjhaBfgWIcnpaqljQqUz38VFMcmwBO1Ql/ZX81EKwdllG/edBcdmEv1B6trTTGE2
kKxQOLpkJQNg2WeJOn1XeXYh7qPqr1qL7IC+URq09X6/H/onfUqCB9komABJzkA/
R0TOYlQMBgsyit1mzhHBGHZS+q1bpkCWWh5aRpBDW9LAUYaR3bttEtN85M7tGnRO
ADkI/wYCZpCPctSJlGvri5PjkY8PFe18wNQXdfruMlo36lHByF2loJFdckaRFXFH
ElPi7PekfioEZ4JAt0aMSfOaAAe+KnIT2BMPHaX2xsOU2CEAmeW4KAyv6ceFM34b
l3m0Ub/eMQkVusWGIx5K7WjLnc+wM8AGZylt8+cu/EuOaCfBAXk/Wj00migfJTDN
4SjcloZA3a0rjE+HyFNYeyYs9dkICT8RssYL5OhetK9nl0U35P0gWjvZR7w8kVqT
sMmqse2BRvfenrnV8tHYacK2cVLU1kuiIyX71ZgKLdAYdjo0Mb5flsrfkl1EoYUb
cOS8dG3UH9gKjuZSrQQ7BK1LmnZxOPG72qTLYa3l/Q0nkdBXAfim0wLr0tPGo/5H
cZhJQZQBX1/1lpO+Zm/piHm+mYtTSj4FShcsgOwbiSArsaf9tnKGznmkWwuuViJ6
IrHx6il54hgEDjWY9MuI9R1P22jIV84IY0CtJxY2VHeuzDmySXmJJpvN/XQcw63l
uRmfJ7dynOjiiQxZHissmfLLDg9ZqSUvKq1j5TGWb8Dn0Nyo4KiqMIuXHiKBDU4R
21V7Lp8RRyuV/EDyFWwAIN9RFYPQYsyl1AGRKOVtyB4rlRsTsGn+yQ6AFayFzW+/
NLyzBw82a3XGUG5SGHRA3RpsXoWZRQL97HZnDRb3kEYD/X55r7uCeBVVv1RREIaS
yOapIJ5Cx1iDnoNl1Y+EIFQuvIV7KY5fMqQlnDaugW+NJVlp6HgUe531ZLVbhRwj
ctqy/bElYOWhoumBvd+YaQnTE+9Nf9RtlK7Rqqczom3iKfSwXIXSY4J4k+l7zACE
vzcIebbvdxfLnXu7WgmXnC+57gwknp7Lf4r5QheslEBS8cdw40EmJsT6bwe7yqpz
zPDAlyJHZ4v+yZh6NSyW9GuFu5Vcls3sTAuU+201BRDG/02mry6a6iVO8RZI00XS
SMAQAHNHL8VTa4dM6HsVm7nrk7ibdntze/B0jJvHsvcWn3zbhvAhDbMFVOh9Q4mh
r9OZyw8uRvzqXxy3sf0bhWdkeD+hMCd1fHrGsFkLpj0flIy6JPbfJymBo0rwtnLU
dNhqRwonSBHx4NdpK9WiOIwMoehrHJ4MHH2qYBocykR1lqXeFpw+hJWHwjhCCKch
6DVEzYUswJc14umiznhRSZ8s8+CvSDheBMepXkznYXI9M7vFl7TyZQi5ypixg0u/
9+i/dntaO20HVRKfNsTl2kZND/b+Ud3uZ+1HzmJgjPhDNPwlasg8gU0+UuDZGZN0
38KGf6CnlnOWqOve+tvdQjTSZYnkLIFOOkRI+GBd/u9a3ivgZKUR/3xYJ3hT0M8a
LnhQI4W0FargcVLJGx/qRa1PtGK7QghJoxnJHGFloACtuVrdf8232ThCBRVi3lN0
xMnBZq3SBHt9jr1nggJUIh0bYxHT1n00+zC1P1rN7Ue85DM2lQAyfsHTn+iTQ2jI
pH9oaSAabzpVvQAykaf+/KsBeywMBNLSkiG+jz4hyOms/fLHr1aeqQpzFtUuBAFN
0JY5qEOBvUonOyGwdqzl9e4+GHiQZ4ESNWKdcCCVmV29FZ0LSPCY/hHnZ2ZI5nH1
5aFDtZTOHply5pHvEy3ktX7rZraIlHmqsiHVBNpJ7ahkycAsDfQC83YiFVyVW7hB
9Ui6jwqca+W6Qfi4ckxQwI4FdiPjKW0kCkZPkGQypEJATWonsTk7u+7w0zeyGYeo
NQ3S6brJyWnPIzGgEdolVhbKsPIgXPUJl9DscJTNjcY1mvRdTyGO+cNP6jczesSD
W7Bse8V9KX1FD4138RtSpm35FckVFicMp7J0Co/1wJY1iu1746GgxU/3Grr9sJUt
ps/AG5Jf85eJwEOZpvgqFeL3mNuAwR7ex7pc0xuj3WwzaR74afrUwIgQxfFqn5RN
blGBomQ2mN8bKXbrNCYnooxi5MQALPBuoEUe50Hoalg0JiFysejwC3ceMHkiM4tI
8UXwyuQG2v0rlltfJQ0WFM7NVIHz/W+hqCFadWrnc6g1b3I2+thie2sq50HUEs1x
LNeV0AiW+zPO0Ra56Fp6w9PlfLgawB1sZzFXG4bY2IQQlXI0/0sLvnu2PGpBby5B
javpxzJm/rAaBt50A/krcDMp2BC107anxZWWDOLqGR2C9XZMHRSF1SGU/De8MPLM
pe21M29Uddh2QVW3YRmNIiBeySp4W2yOYKtZGcC7LQcWW2DsdGE5KMAw2pVJLhz4
d8y6nPAj6IX8yaHAyCBWUgDPYtf5OfeX/Ia7iVHdI8fwQVDqflwiU27LzwEjR5C4
QrWG8FHOobssyYyohIlI5lHVmJS0cupb7vSxEfzQm51J2WkFWu581v9rQ0T2AxMm
NT1L1ipG+mYvGt7sh4EayT/xDFI2C/44lRGXbOL7T/atTUf6MADHs0g/+uO+7LFN
f75jtoyB8qkxThcvpz4MqVVFtv0kGqg8euq4X7Z7YD70ejHtKO/VRvbPvbi4cJhb
2qMpo0o3Cp3FF5cs5QwZlBh15sJxTUWjKISzlig5It+OjC/0uDFbbSUmsyPn4JTq
M4EPXVfskcu/crx36LNv9e2l5X5NJrX7z6jnhlwgtWqrLDtaXohAEj5njnzF0CCS
+zmtZ7PA2SWgpEKuruAMGswnsucQEI9lmYbMqIW+9WzW6FFKNVfcekTux8/8AHPf
hBAXBpZLS+/VDjpi2KaOHhonKLxyau3tu8BGq84soO4uQH+fU7Oij5WoTBR7flVS
zYeyg7V5InrJide1/RqRQ5VquMpLoX7XuGarYURFcvt2iTM6U0L7pq3I7TqWriLD
taXQZFoEoE92dnUJEcVHm2n7l33570VY7aJaSRVRE59bTCKdWHEBPhkg4b+hZuj8
yx2x8C8uwXo1eVrHxzxPoMTwCjigJFk6EyLqcmgbDTqT30xiy7PVqpmyW6X09QDB
qOLId+DwlipN3OaRZG6ps8nZD2g6OCnuQav3DtezKt+uE4sgfRbWtMrrffiYBqRo
22LdeMvJNk0FaIMqZfmStWOphTMpS1lyfsvDYPxsI0MkiOcJWFnoggpkfd6H/WEy
bPsTPKO+UMgjkYcxReVSjosIwoUbkuf7COiBVueijaipVgsiq2KNWmPN4ZO66v/e
2WSlSDh9CfMVnmXl0lvhVZdmJgT54nQnUsU0wyzOA2Tc8nlPfCUmErTNQ7ttuZ1X
vEI6D0Xruoy7Ao4dF6LpeafCVImsTdYnuOj81aTYtNQBBcpA/I2BrOnXyn9lT/hg
GhDKh6sKv/PIGiU1UwIGWaImrWvOfQNNLVNPfix6YED8qaYfFHJSDBDsSoIUX5In
uxTnkiWuQGLEOYZ/vR89fEnhbOoQQlsZSHu0eSRsTC4N4Iugy6/M3XE3xh6LZAoZ
4EmrYmaSZtFp4YsSLMJsGpZpLi21/rHXY3jU+7OjR9CZ+9ML8XLDZc6+dXYaHUxn
OiV6orqOSRUJbhFXxK3KkkSNjoxNIwVrAeVNCEK4kwBWBZouWRTf7BD9uA/AoPv3
CTCn02FxWJq8zHYbxoBkM6Ap0yjTWMaPNfvZGu6gUYdUUTkKKCmXh9GlPBrHJAxe
XW2r5vpJlDElqdQHxQI4RGGc3Fw9OH9pu+GPSkydoAfwvRmqgE7xGPogZjBvKp4F
TXFuUoVf4opK1D1OsWeQbvLNQTvOmUuKvul0WNL39xiFRmkvuaZqWa1HgkL7ns/J
Ix61FwNKZo8OF2inv5ppLos1nymO7HQuGHUmoMjzCf6DuqVluYtCNmIprRkkCmtu
vAtGxevCgdJFwU/Yc4UpkfOm2NdxOD02ZFMUfwbr5SIZj+ifSB9qRsOBBaeBHtfl
bBoMAVDHSmL5iNxqCC6XxP+zhmN9h77eibtJx05mtRmU3n0NQ0XVAAuWtAuhrqJk
js9S4e4UBq5XonijhCLKwENx6+wNL1dQhTIdNB/qnye5XRbzV+u1kLNPqRrqbeMh
fO1FWdTbbvRtxmq6BnCFCB6QF75ITlbMbB0cVpPfYzcGRbXEtB5RPNKsPbsc07kc
4d+fenIuNaaRyhFr9zMgikPrY/ZSEEGKjDCaYe7gi16y3vORDLSio33+Gnl2pHJ8
Q1LEjS19+LW2cXZYOkQY67fT5RGbwNgWmJaBttVvjPHf3n97mrfWCORXviAQsUT0
2R47refvQS4VyxyE61jPjVhbS9MKpWL0nJ3tsZCCvQ0oqN/eqLmjPbqINEmg4+GU
85igAEC2SCOUkAuRsrRYOZWsFXj5iqAAClPMJqUgt6bIcnDk4eIWPnTD8tqXywH9
FK0Kz5n/zbNoTD/mSmwm8vNjNcR35bqpy3lKt7So3OJtD91PWFFrGPRrTnk64F6y
M2v5nAJlXc+EHljjDpvtiezFPZPXGpYffOjujcjSQK/kwzb9z+fCeA8PSSLNT+UG
yfVlBNs4nrfkfy/juAgg3xphYw7C9242Lkha3ZdVWeSVcWnhKtWvv/tbM7s/JwHM
r95sosis3UfH3ZN5cjaoYlmj14A8mBlr40K/87I6aVQJ1lPg4ZG8hNkdQyZ3x5r0
1ghOqlOY0ZG0XqAsM2N6ZXRm6GqHe57epCwIAWogPJd8d/ZJj4e+nV4brwkI6CUJ
FEFtn/ixMYkF7U4g4BcVMdoW0h24El1ccSaTo52nrvp28jJ7pYqa31QsYGBKwBMj
xTjy8wCDkX+h8HN1qZwyptplqzHDtUq69bpAa2LtRIhA+Gc0ixLOI2UZSstmuFEu
zKxh907RObkmI+Rt5zAF+A1d9JtnjdGZxYAAEHfSDPJcWhi2byYxumbEgRNpw3rB
SNemtZo6ff4/Tt92YNJ0WY0An8jw2S5k6HjErm8FzGungQH51Jz/LzeRQYqa36Ar
uDF6nxX4hr8sg4ov/12rUgOYvPghDiKq+4cC4Z6ucpQStToV/pCpM0OTFCg7L8Qp
dvQ6TbG7iwmfnv1aK7ZvjFtezLw+h45vlF2oOjAtA0eLhiUD+9UWjXCwppeZ5PdP
1RcXo56U3oYyklUoHQQVUnOU3TtiFnaecds0/uFY7m/jCPWFjmQz6+8S/ODCCm0w
/+59nsAUOSXpDTtvX/7Cw9QYNEhkfA7lZt9D9E7fN/heg3DJov/6mJQvc1rl0dYi
Jqpf2NRqTHkazjUS9ABgfZpbMV9O6d0n71psqBMpZZCizefCcLU/+VwnPaicOV1H
XN1hYzN6UrTEnK9Q/6JdFtDbCaNam/NzRlDADF0PUMA+cfSDikt43JcJBPCFj6G9
yLE2isuSfcz5On/wdzopjF/xfqwpeC1ftr1PWhyNUHDTNKRv4XyDWgo8iWCOcDSi
aRqCQ29i+PFLsz5GZ7RSAVsQf10HLtU6P4Jv+8KlDgkrfAImEPD5enua1MPDkp3L
jFu4ycggxm1FO4D399khW6+nK050D8mSOQxWTgmUXMXTyoIdLgVyUTtRgT8CHOkB
27X1JjztwVJ7dgWWW58yz6UnL+tRbouesQ7KLjlFT6iYMunY3CQ+g+lmjdIs8CfN
xVmuU362y63ETMvfc4osWSkS+IAt68/4SY9K52D85CUmO6fQNteF6GnsO7KSZ+3X
vQJ7UILrPduaKtd1pQRMxXA2MveWriltVt7AlkQ7n8Ey0EiMRLIBYcBxu9vmzUEM
oeF+B57c0BI2CJoH/Js+MT96UQu23nLACxokrJEL6HAyhFXzui5/NZGgIjioK1n6
aQAeKPPZ+4nXcXF68Rueck/LP0hxwZlwjk1C8zct/67Lhe4Xrn086V5mg8q2Bb+0
nPZX95C7D/HU1xqnLQAmd8DsNYVXMDxt7wwaIC9zN5VB7zbGFygr0Od1M7WOVNvN
QmjGKOMW7jpWR+zELbCaog9Hipl/TjddSfy31Yg78D8OtzUupUXWI1FfXtx8jc7C
+hMXWrb52vYeLdUGOzOoN165W0Oq8bB9ejGgEkXSuLYCrfTYLmqND/DKuCw4MBmy
0GA7YTq5IVYzPWpXA3dDa59RyTbw8B+WsOeCDQOsoKfy5VdkQvaSO+e4rBdCULg9
uCn1JchEO+lEkghJzE9jJWLdOekNfS2eLytesvZo0BWN2mTULpyyfA9uhMIZryiH
9f2cW37pOH/TOR4/DtWLP8foi4ODlmpSI7Sd+E2j2Bo8RlTEqQY4tTd+C1miSo9q
UH6xdCrzJwlmsuP3fPMYBdieyNZKRJHuw4Z4hLOveqc6jL+XkCqfqBabo1c2IGU6
0qUSVXt8p+pASRHchDGjmiA+GviI8HuS7QkLO56C+uoViuhOWyC1/te0iLnmdGb5
czeoGnsExaGF1jJZgPXcXQN3w2zlBLG+fZ/PjGZuAhnxElZyksnmSg3ro75U9xua
GikJMRXeP7hErjyCeS9EuU4m2LCAomyVGgkIDThizJcT2rNKtrJcTSenOl3GtHC5
ubsnAM9rXI5CMlYU4Oo+oKaKVtNw8gHK9871YYmCIVEo/3ex8QU7kq2bPvC/fdqt
SmPkZvy1IPR001k9ttYxMkFvWHvyWNtg1OPrTbgG+/1AZMyJ6k/jQ4iszH5A8xG/
opZndj6eFRjYCLKjBOOAuL3M7RV7Ab7WKmg+57Ki1hVMVtK9TQsymvBQaZhpr8wL
tywfx4tiQbX0Lecp6yKzHCPboyYeoUTJ4sftlHJTTzsc+zKPON5SjL63j7dOMWwg
l+P03L/4irm5Nts+4XJ3E5s/3p0GktfGO0V0gR4y685PBGZCsGvrq3FAJnuB3SbE
RsiGkySidw/iIjJiAdAUUTdBC2tXVnubz1W6Uzt8wE0M2PTFuwhDpNGpolPeQRtW
b6qH5ysdcJLCfQy9aTnK2wWtVX4JlX2P9CN3RrA3h9gWHj+U/uTLJpYGRfTdaHGj
KmB+fdUPPbawudhIGt1AddeqIO0kWUy15cNADl1kQuVNDkDRd6hAmgHfxEIPKRFH
TvWbsBpc34k6+BzIzO9dFJHuVNxNikwDweNRDhpwpXAA3O+cFZnINz7xQuNw9/3u
GQgLPHpa9oL+XiDspkQMeT7vHbG6D79DAH7l8Gkt0hyZ/UUCVokEbc0nDDC2p/lI
AeUcZC/Vd2sze54HVgOSsrZPHjN7xr7biHcMmrZ7cnYPUyopuv4YqQdfy7XgN1DM
yjsDlfnps0tvS4Sg/B5Q658qbL9yQGaFluBMCTzxKi+4vuaZPYdaqIDotzeMtqDN
3zw4XsFEb7uOdfgCDdrP7aa7hjIPGFx/Gu/3/5HJQeWRMpTd1eXqkCaEZLCGi+RA
HTTlOd1vsphv+CnAqOLCqyZNjSzns+82CHnniS+0hAyLIAZDtCffvyUpXha4N8x1
URkXHqj5bJrNJqSbROLqMY3NpV8hFyjuQ742vm3JVB+EnMx7vdS1bbVzUtoRgPAq
OJsGNGl8kBOfyRvCDghN8vm19LWmuODEPtqFtvVXXfM+zn5H/xLhIbCa6fDGzGlY
RveqCXcMEjKZKnC2idE83yYxaDsXM+8Y5bQs8fbEWI1Q0cjzkNP6DCnP7WrbCaso
iRDswjYnIIEbL1bH2Tk7YH/3G1mAjEIeJnhIeaC6v9fksUKF1BL63dmrZ2jc8Q+G
ToA8J7G7Gf6G9Ht0dfSa2oENZcvLtLnGOKBtLqFlT/uMazRyjHGokCVERI47mR9P
55nwIfl2ZrXKBXcCuiEZsusayUyhMfsT8BE4P/z65++2W+V1b/ncY4QfYR++04OL
MF/YElyIMF0AD23bk21Jeq1kcJlYQ2s/Jl68XUP6KkwVi8UlQBO7fw4PEfjYP3ME
b4OD5EtkaMgRZEPH5HPslk5cDmUo2nWEgOXhZJJbPWPObjR4SAUSDKtxxlfa7FBg
VffNF3d6SsFvqu/8dPRA3ynPo4k4S9o5gBLw3ScVSalNtP/WwN9JEB+VJ4+ac2io
a5aalpPlKTmWW0vZnUOX1e4pAru9ObcWkmaEsKlEnXsv87pVBnlYiuFgaz8S1hi3
0IhpMAsMtG3HHDvijhVlBNy/H05agsr0yzYYsvpgXNfrim7lx+wwnVhsE+PACc8W
p5yUahr8Pw2l7FQVlrH+EY0lW8lsXMvFfOlnwP0Cq+EczhLIMAsXXyOTEn+6l7dE
ZYIwfH6vuUiRA7GnAf/pQXD3rDZVSfjL8C7LFOf4SD9cEDTU5WYG00WIPiYLVMmW
xqnElshNWAbU7H6XSemdegJScY97IJAKJS7UCgF6/X4UT3TzkV6MOu1vAvZNRgYc
cCoEhmJPSbzOyalp30RXjKWNTWz1WFPWkfanNblQAVeuTLqUrkR+6EtaSItwRxEp
uSAFw8nMOEoVayr6BLcjApBmoE0ZE7p8V5CXHEtN7JR6MNSYljrX9izfG37n343f
OuL/+nUeG7bWOqXLxmXi0zuH0S1uFwm/ooKfeL3D2rLxJf1yGWLcaJaINVqgFbGi
1Va9kP1Rm1r+eusVwqlbmJzaNDFPX8aqgefEmbqx/MDjxrYPTh9G8RysgjbGue4X
GOWzJY/TDOQ7XCIZpq32Os4YAnO0iG36yvOkX7ixN42dtUy5kvDb3JaDYIMJe1ik
C9dUNlyMPD79gHCpipFENaDD8ktLKBxLgODdmAzXm7qK881gZpPF6tA45Tm9l/0U
cODLaU8heiXExnHaVTMaHnvm7jgbh2mxo19EGJYP2a78EsNKMXD92St65MMke6HA
Sh8DQ8WVKzMj2hOcZ19H9/8SuhPMT73yKxgcRwWImZKLo9DG8PgsZXH6frPXrjUj
4KLd1pYibMoaRkZPY8QTkz7VYZ8CibdSZZazVOmBPnsnaRliedMHPt/p7YGJi2d5
gksjVQJYI6kfuVRPWGQE70QT/sJPUN7N4WAI7vHF4pGaoy6MsuuZhFXNeBoJexd1
cUQBUNt4sDORQyXMR9z6xyyiWlrxVdcsBlaqUMEZ4p6ngltiG39z4C3d6hgSlSd2
X8FsCpc5nBpKIMb+qnR4rwLm7E+IrGjypFGNvT1viN872zRGoR2hTzoQ1q0TIUD8
/dLMM40DGUrZdHH4yg503wcZGoHR7hdLLZPnozTW/Wg6InAcO3z4Om5HbroqcOvi
NBIS8VOx/Rot4Lycz4mb7mSkjsH535W0VF+4wuEZty93pcP70hi9rFRXx7IEEaIF
cD9yBX1gdyoj/reURxsxE6vppXwIFiIlxpwFvyIThAoVvM9I0iB7anWXBTMrXv1d
+fCFnKvYvucApZqBpe92p/60fSuaoeMKEVmZkV8vZMXg0E+wWzAtD0G+0Iqa8vlz
ICMGukScJ+e6yrWuW1CfxJB0x3TooMolDUHRSda3Jqz+afEZ5bBJ8VC8dWcgazvV
RzagR33feoZTVczjJ4v63R4i86FzfWhwdUcr40ioXkTWAbu6zlvqYJIGCqkc8gg3
rcK4e6gkRbbL9+jBGB1ZtorkZvGiXeeK46tqzLKixdN3xowFixumqKHyM0dep62W
NUHj/rg62YHpIg+EPFwiPcPbqYpWKz10h2D0J4UGpfMznQyTNZFMJtVIomWZJ4HB
bfZyxOG6ZVcWZkk/+0mMPNXdaGTiF/5IyQTd0IfmQLglo5JRo6Z8y0yAkEtIWAIb
5qO8SxeHMduDg7Axkg8ekR9AEBngmSL90J1vgbLjPfMbmyW1fZvTVyVe9NkmIPzv
+79ck7yGEDSNZTWFn8LUgjHU+BTgAoIsjdnnkQRObO8VOVBbeTK0zXH2+A1PhoGb
l+NYCtuzJEJWL330v8Z2xSzCFif6urwgFhDLTnWmL3HLT+J+7W8vqn36RHeV8uC5
zMT/h8xkCva4Uyv8AOQ7OrgW7wEbsdgSI0UwI5nnlQ7XUn9umDb13bL4cSFakll3
9Ijcwj+xDiiLcFZ7QRr6gfL0De9L+Z/WdJ0TkiD0I5i6vrSMqKXCdMvOOHHf3wHi
iKuiFlTnKlEaONqP7ZpBJDy5OMdy3pIB+rnypG59D84lEdflzyUeyRawS0k5AzFf
AwJO9eP/wHxa3+4UEnE8hDwytiQo7yy1ELWESoqpz6HFjdcwKm3kWykJqfUcy1VI
sRC6YPhgWvYzRQkJDr5OHEVweWDBZevcNuws5KDae8q0YLc32ESVCkKcM91S84dl
rG3+1N2Fu22hfu7mTDI9bYPlNJQNr96ybiP7r/bWUkTPO1ytmEju775GnsOpK2tf
QVYWiRf4hq60kvr9fDlCEfUJoQP+PUyx0PRBZJ35cBkN4uRkzJBG4kC3ATj7TeZU
qf23PxeLGcFsoj+H3ss9GyLfJUhFkg1NKKZgh+PET9uev7hix7KxXCQAPWN92emm
av7hedaftN7JO6BtecKznOC+ctCcB3Lv/EbM/j0EQ1fteeC7TBTxktDMUho67Qqa
CQ7WCFoCkw1gJEM73AJtq9TpP+XIqDs0MFSb8TglxoZG9wUTlssh2xf4JSlDZVzk
ICimL9wMq8CNSG+ZQF3PqiruzrFlpmQU62oaxQkpuCyHnByKwx+Ba2OpQR3XOjta
lKQjm9fIOMX4MSQ+CttJbNx1foIVAncb45r3jdemtUIp1wAdKU0NupvNTJwZ/LZE
X2oXD4HJn86g7etwInf3kqAqIqN7cwtoDHT2Y7Xjr8sscvpjQnaRzw5yyRvv1cqA
DvItjptqdxIp4kKLQUCtqhoyoPimo5B0EtHETHknSrXbFgHVXBP7FtAPVIw+wcj2
A9O3Qf3IYD4OtcaMbgZkuPxkhmUpwY7w/0fUf80ep4HWCzxMWl2N+K+TuO9SvYfH
JUec6sWZ/N225B+PIu2TJzwg412/e1YmH+Xq5te8xXqTaEtA71iMoTOkG1JaILCj
dyBJq1APIDhph9hjGt9VUP6Sbzz1lgsafmIH19vsYW7M+sY0b+SISHpfIb9d69Na
KKk7tUgxIJ0Oz2GKXHYUVFhBCJ1j/uWZAaoj0Mng7/51hppwUjL3WZCIJAJ7zNrj
L+qp4YI68Olex+zTR6c9kanb3oi5Tw/PegsGkj3ylxG2jRHSJZy0GVNZ/jCSgp9v
NuARQ10r7TqtnN8b3VLj/bs9VNneDpjyjI4GrvkmMPdHw5CRCX8WUKx5yqjfwqKn
HoMIqay4shf9nrNBB/xVJb5xtAdxGRAG61HrMGUEEy2alvz8v4tLnj0b4CTn2wi9
`pragma protect end_protected
