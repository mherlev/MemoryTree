// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:54 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
o5Qy0BUIhm0rDwdPyEz+oUcGlNzVjb0wgfnJKj96Xjvk8LSPtEI3OZee3POqbmch
5Qt/N/zgWlphai5HKxOqpzxgAsMSnLpTm5JDkbnanMsccJwrkeadjzoTv6hvlui8
W6zfzVF3iSvE9aHZNsGKmhMEyby289HmrYjI155Cjas=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 36560)
fAUtnVBKLDsXRVPTu8+fJoU/1GVNKDZf66WYfhn4gKy0wLbbi66hnRLQ+rZDDMvt
gFvBfQP1LzbrRnqfDGTVDzihENttkuncg3lrZpX3Vi0TZA/SSS+HQr3rn6IC1vD1
9e/OwU5iwaKpMID5yw4iOoddupIjmhHxEOfm6DwaR4SE/j9sWJHlgKoqGKObXpTH
X6RX6l29D6hw82CC+RWYqgHtK7KCbxTozpiCyl1Yyuv8DRlEyCpCM7bYofsSME51
Vnvz7MEJCp4nPyik1JeO8Zlq2d3Lf5+PMdV1Xcb5/+N1Pxt/fUeHlZAWH36TOZ9e
dNlUAcrkI9skV7QkKJ1/TFjWZu9zh4nIxvM9Rg13SGVOTz4yJqPh+v+UHdRHD4zA
3suEcJWf2MEkiJ9laUhvsDt9qPIyz4G29GT+/mTbaCqVBh7ZK5Ce/pBTy7RPZUPO
gJo4xHwjKUnEtMeZ+GxkIRn5dXmMgHweVA3py33Yh7d5HRVCnvsc1fzkCGALEPdr
4Ax5B1ZUTCi8/4KL95Q8Z1cMFQjLuDtgXzhDeQAXID7dWPxl71PAnKSMJxsC76ag
Vl2M1VA57Sk5T9d7LtzJu75gMZ3J7a7y2HT1twGYpPPy9YT2F6kCPQIxEIlCyYN3
7BUTPbg2lpIKXGV/zuZD0TM3Vrpb4tqF8ZWnhVL62heGQj7k+0eGhysyzbuEUmtF
GtJCF4JexQH1HgrsnW6It7EY2L7Jl/KLu6yRJnc4lofGYl/+4ow/G5TibF/WjNR3
UyrIlKcVvMGNGotnNBFMRXWpAd524prVA3rMOqn5bs7X8dhYV38lHhJr//NF8uV5
yD4V73MQ6YILwKavcLH2D7HMT36AvF7TcaNcLNZuyTRGjj2uCXAZuk0iVUcKbTUK
ZQJr34ENqliuSGahIUmDogV+gdx2vr6guJ61u3MPEarDK1EHm2Z+pXePX6CBVKKd
QA7l/CCfPeJE3g4E6C8rne5aXxxxpULqZ1aTnpLEtlqbF6mweq9PIvXpyEBBGaF8
PQwMadwI+kEsM4SlUcNW3Uub/NX1ZE1Nssmvxhwqv4egv9ko+rPTQNP5WSvjO5Z4
4XEmv17ZV0+ILjxfoKtowfLjdMYIV11JDt3dc/8jjuAW/j1oQCH+G/nD9vZYqN2U
lYivGCMpKiKnnktOL3UupjLYZoCx4nvjIRnjZTtyHxkpCeqv+faY2mqnAuEN4xY5
BzsC5LtvLKdUYV8/U/f4OZ4OHMabLcF9baQTSTe6zhcwzyL9c2t7pUV6KCFsYQbq
Arq6a9ZscfCNd26/ray+XSMkU6TLk240lg+T3ZsP5jvFPzpA4jt1LC5sqs3MEz1L
87PeNMGv4nFR2isocgUK6w/mE7fknm7uW/bANdJ6Kw/SayxArkeO6TaVlutuBNAi
3aqRnVspHWga04n4nwouvD2J4aPCYTKxRhJn6TRA5Tl7oHgRug0P1pvtVTZX/6nD
6Y3aupwAP8ytRhdd1L4CzO+Zp7u05ilAI3VUBN/DnUb4QxmfV1ox3NnSjJxqOUV0
G6JlWmUq2KxuTu8dtX0oGz9SEWs2wJq9+ZAAZ/u5TmOxbBGNV87nkJQj94iE7K8M
LsMaxBuJJnuOO6Yvj0haKlSq7exdrkxcFWIREAe+Ft+hJ9SGaQxAKrX5lWLQg/OB
IGXsWi7FEshu7g1N7/9b7+xPJooN06M0290Pl/Z3TMETbkI8ThBJW0KyjGckQX7n
tgJAxeSwZcW4ovIe1IERQbM0KZRIoEwsUiGtKA9xX210FZEEFNXoK42kjZJrpgTa
rTSbuivJOTemVpw0j0uOt5DD4NpQ31sXNUoPV4bJ0JQAXcxNxNxPnYp95+ORebrH
HMKG0VAybKKi7lT7wrxqrX35b4fJ9BtlpFedPtS4N6WWiYIRkveEmVqEn/HRv93L
cFAZxya9Xb8PkHppdn7vCKrEtwoiljkqfCJWginM2byseL2lQaIHXXiPPpCIOsBI
biY1S5iDCBR1ARXO3qJaIGdkRoO2qKWhcNof4d2wRLObKBClAKQJa0rMOSVXHqB4
bZ4AQR+UzAUmMVHJR4VYUI1U2a807kGr/dUyV2Ff4Z2/B3YeLuLSgp/AiQApr1lk
H2RejQNzSX5bEp8NuZRl4WqW3lqkOk+eHv15l2c8ctweHbD4asleuT0J63djsFpz
fpbCHz52uTMh8sZnffXiMairKlewbQEfXUOTFZNx1o8EUOPOuX7u43Sv8pFCG9+m
ZUVuplbhgLVgE129GDRc/zhFvbt/0+l8Goc9le3CbjWn52U0JTQH+uUWvCwpOrC/
IAG3dWZxZvk38rr06StK8QgQhdV1l1gPUk0teNCRYxeh/6unth0sZ0qY7UTw5gcA
eJVV8sNzyH6XJSi1uIN4pcxPstn7f4zIby4y0GaGzIm3xZidroHgjd1AyDPKzBd8
Rks6wswP0Mu57Io9RrBjiA1lFbJqZH9F67qP2HNmi4Uf/wkqyGHF7MjvDi0vrsHj
chW2CgyhRCa1aK6MFyRQjcux0CxTWGBjRIP2lUGnSOplHwsFBAeYtIXP9yr3uBYI
xoz09dxnt40lrDr1FfQ5yHbL0YbT3q16FszC2O94Y52eVoSAwDb2r/ISy1tTY6L9
HchedQhBcLNS+wYKgNL3eXR9YZSkuASfDW6RU3bYJY2R6UEfnS/DFi8R5rkMnrsK
ys7YRgx2bdLRXrnOM/n+TI64Nh0TK1feMkO+tGEkI+fFtgmTjm3NUOtANtlpVqvS
iE1VL43RToNZpWhNmnurhA3/lK/ZXGpiQcV32NRTCuSzed0bRAs2ukCI4/BG0rCb
4rfV/9/AmlhwEQUbPyYO4vziqEeoH/9qS5+J6V01eB5Cz3NIAtcEuxZCQf5D8X6L
yzaDZEUUSNvmgIJHgnBAcktj34LVPqMvMK5IzcFJZ+Rv0fw0aE875JNcjMPESGKz
4yQg0BnMp5DepjlIY92BHizadiWSgmjUI2wBwA35wJ/4x6m67k2aBMA0q7G8sqxc
28ClwDMN6xL4ixtlX7jqw+ohjLKXKI5jzUfe8OyTY6gZl7SqHo1xYFktmIy25ima
eGg7x9cT+ET02O7cvZtwUDwhxBCCN67/vJ4DBAhwDWiAc1p5bdK+BUNeW36HyTOZ
76ATODHIoevIE7npbniO8u4C0SacqR1g/NdiepLcleO/pAuC6Xif/GAvRYD+TotE
gIYpCNQ86LbX5xdo1vWtBv4HiBIAfqf9+WludCx04n1a9BEpEaBi0f3Oel1mOTpH
fBJT9E/Bxvyj0vkfPc0UxyWK06YXnY4jnsQ/0Mw0DuFPtpTy8vgh25J2mU2V097e
Qt22P2imd9xKjiVwmZyXfm39fgan8/YyVA7kvJ3fCT3atqQYLAjLwIp6ui3/fVR0
6j9gKOwcIWUL19HFP5GsmbjAU96Gxp9VUV2hbp4wvd5VYm+/q/bUY0N8rQg9Xwop
zn7fk77XtB0nsRNoPX2wGcUDZ0M72QWmcXXRZeBYiqwxBni/Z0VQu8QZalDaqZnE
1VY9i6GbEp6wfchdw+CT7U7hSBi3HL16/n3aZE2AUY2RX6cxrpsK8U0FqQwFh493
93JjuduHeZkMSTA3mH55zdmGiNTpBd3e3+UYs4DqD7sOVlw6obfq7o8KJqR46PNb
l+vlnlfzIINJ940JVDUHc4TLX/icaTKHBBXKtZEFEqdP3M5pAOG67Bpp+9ByWaQ9
10T/5w3zt9Yum/rIztrxngEwwEo2QsReuLLKLUyb0eZoLc0QwhaUOLDf/54BTCge
OdFTEUsF5kegwt++CaXDsvi57wXshGgSuax6hDl0TZxnS0I2/aBgpMZOdW6hCjA8
/cYLIH7fTT2DsCSHqrOt4bF7jQhr8JUZrEmp3uG3XXwGO4Oz1lgOZjzVORNGJ6mP
2iK/8Kh3YxJLcMP/6gLaZ1vR23kp7VLmcxnCUfhxQwAxWCnvXRp0QJFYncFEGlkD
hQr3ZQ3fxPeM0X98pNrKo9icgoNxW1bU86TqlxnSwvsIRsRYzi1b+HE/xtU5xi5d
4NNlmHfyr/TEUC2vjvw2KeLUneDdKlt7B9lMciHpXMwcNmcT7o8BrVCxV0PchSgE
pLezTmGNVEA8MrMn+cbRzP9VvOxqV/Mv9+XcQHNIqWT7kfbW+A7lKJVRo6ORLPbA
yAezrDXV2/QZ0KoG74a67/E5tKJ/c3koqp6xN2VvEk9OJbjG9Y0x62ev419aK4l7
RVhSoJPHUCBqkPwLh+a2JAaY4tKGxGhCay74AZ3N1EAsGOsmm3j1EjefMT+a6X2G
b3UNsKB/qLZ4n/0G8M/CyAHlauvvxKKt58rY/rls2Zu1LK1DTMUMciGJo0v5yidY
Um1NJnU3kIjGRkKlisd6pS4lTpDtRc0qH4T/bdtcCTCzlTn4k5hp4uf/8TzevXro
AvcGvmvVwaAa16cKk6cuGbmJg5M+27B7D97/UN5F08GeGGlQXxXVK1LDs/WmhKeO
JkEsrwsLWwSe4KV6pxontWbBTvRt5MLQqknOZwnm+oxw28OLzMuowdj1yzdE5i1a
hyWgCWYykFKKconhp0iFlmCqXMAjYdoKBsNzxHMGf9jC5ECu5YtJOrP3c7Er8ZxM
1alz+N5G9ZNrh0lWo0GPBkQU1E59DBZkK06Yz/HztkbcKGerFELDjcsnCH3FF7qw
7SWSwv2u5i0Xo12awbd5T/CHVgtA2IZUBezvyU6S/N+GS7TYSnnnbN8YI+DNwK+s
Qns+FD8aS5XvAL9xAZXLdIRYX9HhXNe6BZmObyNcRI/JhgGJrB4W7L1P7YkSwFy6
Ph2NlZdWEEqJcsWNsQOsNIDCvu8wxQ239qAbQYq+8byqim+KwypMRmrQqJ3OcIMv
vRp1A08id8loypxu5kNVUf/AdPUU+cVMMvmytIvoza+Uwy6QoMLvusyR8HHrKZCg
WNfRPkHHdNOw4rC1e0IYP1xKAk2JCKbRBFCA+HgxtHV5+ZJMSTzgTWCx30dpt9Fq
eYOyXEeDCH0mI+fGvsJ9/bTPRgNSVi+TmrGjY1ZhhXqLLemGZAuHmGv5T6Pxrt09
RLuN7i9ahL4jZ1GZ8srTlVjEL/fAiurNa3ox6DMcoEU6XpaOjf3FqZBDbatRK0wg
FzefaPg2nofCvviTs+8E/x4+O+FTRwangSFOtUmTY+7fxdubaL9/oodIk876lHrM
4n6WGPSOqlvq2mdZiqkYXUc2FwNrHtp0g/zc5iUzOAAUR2Slw3UGx/gguQ0gLLZ6
si0L7QJ4CGiXTDQv4OMIHcKCuJy/DCJLtbhggh/IlfbQgI0abJyzYpuMeYUQgvpS
1pL9OS26GIFymhJp+UREWGiJMSb8XzGcYt9DE5H7IToHYwON+0uoBzjmKnjbnwsS
XmFbOts/OV/gJLBoZzIOYwj3g6pJ0Pi+mxX52xve09RXmajLdcp2DQJdOcPu+8zt
1bCorqAr9RcpgXWD1cMZ/jlsaQcuXFTBdq1uFGfmE48pHO4On5gasszMIh2X0OJZ
YXYD+HYTO/lDHaVFE8oKg54GRwLIqNr3lXaoPmQ5J/qkYs8KQosxJtxyofF20r+1
c7ija+9WWgtDrELo+GMW+v99W5LC8eGodyFXlP2x4UqUaMatiI1CZg/SeUyd5HHp
sPIfb6IXA3ZNlDyQEblCwES4ki3fj8k7afGyWjljfIcpzXeBZYvFoaB9Pi9agrbx
+KMILqyPr/LTHgytmkW1naknNxCUxqeZL0bjjX2faXvp7wSqncgEtueJs/3sCSLg
XtBox+rX6EGVBj74NaDhWdcYTb3BSosKh4o4bYmBbBANzNWZrvunyEI3MxqwfIxR
PTQ8L8ARIvNjxVMQc1g8uWw+T2pMVcM/fo8wdqkppgz0rm4b2T+hgGb1aEtEjs5/
6NJTi74D+57sTwDKw+FIGtGDsEExlzknoqeU2xcK0YI+bmVcVdIrCPJ8/Xjip447
PeEEjoynMuV+v1ahbzjMeHUJYSFObph8oNi/mua0WvZHvC5ecWCsSQUBNvoNwNK4
3EMUbJYcfuqgf5kOQ1bTjp0E62V6nytqaIc34fl77NlCFQzwBDR1DVTGLO8CDdAg
TqZmVtnoFKa0Zoe9/ekvr8C/01oHnQUfhPwH2kSr5qDKYVZeSVZ98Q+4GcdHZL1I
MOKUUrtGugdFSeptS7B56WdJcwwcOAOedNwMZzDzCRHuoJdf949mUvG2lhYXpcXj
fKEFQpITjnG5/cB3R4S496+X7qghzc7xZt3X4LlCIRt4H4FsJr2YhUkbVyhDhK8B
QrD+5Kq+pyMmyR+t8mqR9Y5upUyh5a2nIrDLObIFdWCLoxVAAFjznPgX78BO6s6D
25rygQRAvMbaTROgs7a3vabqZumkKdo8lw67VoKiGLsy+nwpQPQKnDoOpVMwDEJR
Dru+jotiB+OP5Vdy9VxRATTGToPts0/QusDq4aysImZswJfQZlvqUtabwoJYGzkH
xXyoOWyJ5+sApqEJ83ay/Ca1F3vdXLVbDRM9NJm6/YCJD/3tpMMiw50pS07xBotn
D13reroHxGnDNkBJefiKDBnwpkpEeo/l8j8WsSMFhobBBz7+wBvAniNSoFz+V/Sy
/FXj2zU/u0/nTULleUWNXwX5MbqpEISfvERXEkq/NydaXj0ZaJkcookVVJoFs2Dt
KiJAvKI4nrFNN4WNm/Ktd2iyzCWOO9RRn2oyG+msOPGJPlMh6qZpLua0XsMfBvan
D8neP7iuwXmEf8Rbc3leyiz9aqHJ8SxWct391ZMDLpz0qOhTSpA75IsofVMxfjGT
7DkY49DzVW7X/jkMcvHvVqNtaFN2ZyC5j4lcJ0MFCi4ilvj9i7L2xm1ncakdYlDM
xfKXheLNBTPmFjxmfy7cN4R8gHop+0/C3SbDvC8oeyjOVxz1kK0QmLm3LFapopxM
p3BgdqyjRcTmCpw1Kpn0VMQZTxhsVzipbx7tg50UYcNslrm50UrowPW56RaKWPMQ
CNucCxa227bMQCkNZtPiI1cRYjmUBxWYueU0e0vwyXaf26bAYjlMcU8szQGipuhi
EbTJnRGkg6Tjw+BxYh1iQoD0voYTvQx3ql9a8Lm3RVz2WW7LHVb++IEXIndscMxS
hcP5/tZc6qcbRlRPaKlroi48FEck9VQri9mYGr+6dCZYySHLHrI4tNsBM/qZ/x+d
/g0Ng6jLyjszl3bFB+JJ4Xd74HuSsMe7BDc9KaUokT+r5CSe7a8W/9zTf1mZ6v30
Odib5isZLMXhqBxs3tMyATjUjLuEe4SbuzvqX34ZS2rVWmRjtTO5Ugl01edCQiHP
qm1j1CvxOyy1N5Oq8xxQhsjrtGB7jZBgpT8LBwK1eiICFrCvt/qZMJrjpmjcMu0b
1ehEWjti/EahYUSp06mgrbY4pZ6Cfx7galL9XgCOpmJSJFtHwViwvwhuOlgbKX2u
Bc3BegCBC8WaSNMYxJjVpATdv5gFDCksAQcVl2Sre51KUZXmFy+AJbpgGAlXUDc5
yxPXG7XrZfsX4MPHHJIZZuL6v2fJNxhJFViWnRjDQVA05wNT46Lk1xyBMC5CC2du
EiwnDa+jjPiFwC2GEDWcMzdh0ag2blwgzYJW2nLBkOC5M3zkGB88DfXZsWxqFKjh
XDVUzU/5I+ZnLKk+lIfvT6k/JPAq7AErfMVoAOHXz0NAkD95hzegrL4I/SCG6T4r
OQ77Vj6pHp4RQtBv1jeOyO5H9QpWyVYu9L6lEo405oSACL9+QwGQ468KQKdzLC3A
RXNs+X16wTDRDTHGQmIBgtN8kTGZFdGhGDwGcB4HSO21cHDkQEw1yOJwQD/r+wev
Dn4YbLGQDAs9ytaf82ygQY5i5SrzTQKbUBEOUsDc2gr0Coywa21qcOY7CEl4wREa
A8RrsL9hwth+E6B7bdsroRWDmL1vhSCFDEo4swPR/z6IbvcM0wvYGlXaConvqtgy
ebnkOjksdk7HYBFukjVeMEAFykvuuW2MkRbTPmJvzUsVMc7fwWvBSPftHgGZL6ro
R8GNqZHDLeBSKiiKbd3KgIqF15CAK7v066IkeNPXHDqW20RKkgaq4y+0CfkH8Fsk
uHQDMYBo+QmvqhYb5JDXUn/+y43PI9AADJt62qRN1B0LaDTtE4K8cVDuP2aZ8vYY
2tzIngmJvw0lMLBXstwoNGRLFqkxeLDv4gQhFofWs5Me9ltQRdnW4Q2LAFvCOwkx
mA9tvDmaDuM8rUxY8Yq6BDLH8LcIemTbTUsMBAly+OwSr4iSqL7vLmDoDSTy+vtQ
ZKILQ2N3662+7OP2mq9MFgWeqj7rGU6HpxzOUFv8uSInXHGNGejEIqm0hlRQPctt
o2EH8+OjNOSG27ptDKbFR9+ArrzGJUcKheb1qDwPgAJeebKRk6Ul6PACfv2oVf1C
txMAvQwI0Zd4Imm9XqnXpXPrN88VilX4S4uijPaF1wavp0n50ZE90hVTeuwamfDm
bbkMo/lCBOr21Pq/iZpeOo+ZyXMPCprxBtDg50ArBDx4f6LmLVbC9WsJi2sBrgpU
IpAyORfXiJnGgqJudWzlGQT+8QREoiRfbhvqvYja4o937u0EBhn+jIHN6ggomnsN
f7twjLM/hAuH5H7ZdcFoHxW1Q30rC3BEL3COMfUThdEQ422aaoVqH4xYXPPzE7A6
45wPIbZSiwX/zpAOvK2UxXUOHWWvGrLs1JqQcc4IucpPEptk9nYUbFcmxAo6ZUlm
0PA/Ud+pv7wiLmBlqCAdmCxhRlOYbZTyaMQ7zShXFY/tD/MHvsRcEl4LbH0Gfybe
uCQaMGzUjC1+j1HL15HqXoENXesBE5GGAFiir/lftiNO5EaKAGkyMarZ9QSVULNR
i+0hSC7H+ND+FpCrVWx1MURjd8bBSoSGIIt8oABSA7mDMG/17mxzDdVlycatXhEb
2eCnaqXrcvxlS0F92T0WQvkdR4HwOYcpKDSqv4WkRCf07E8JSy4Pnf+S2YI2T7yD
DYfWeMpDiyYG5jZBMU0e/TUCu9OYCEz5W0rtNhxndB2MPv7AZ9ibvXhs/DoFmALj
coSrfo2af6BYIzbFy5t3tFFpYcxarMOYSvDOwYgbjQp6VX7yPZR/C81grYinek9T
io2LTj8e0djfHoVXZgquOv5ve0nSoJRMy4qCkHeHGnfMWW2TjG2CYf8RGcGv+ylP
7WkO0EK2w15X+R/wNaJNBzLQWX7yqokBj9WXfw6D/OhNmrrZO2KnblaGg38G1bng
n1w4VCyljah8GohXrvLBfdPTIGrAShgmAAk6CU3a0YG+ICvmPKp8PiGD8/7/j4Un
29A921yThIQHu1ocD9iF8sQqqLwDCRBkLLt9s9staodqX36gWC0vGD4D9eH/CXvK
Qk9xGLrJktJS3mrO+Ol+zaX+Fla9TYdWEitRVo42+fIelENYtwMjLML8PC91bFa+
Vu6AKBFw2FlNaSFBK6gq7SBKMDjYvoXRGaDoS2nUoQn4WI6LhCP32+O1v3otI9SA
PP9qecWUjQyUE2f0R1/O/D6O9tvJwk/XplqTvhKA3JV+qjJhTtpWvUmiE4oSWe90
0Mm4cuH/HW5jBKMk/twCZ4DYfH9daUK9hoPDkAJgCqfsU0s1lzQjzDBPrafI6BQx
yqWgj5GGahHuVECPUtIyvTa0F9+oudKbdknX5R7s98+GfJkRgYT6AFXXLU99plwP
M74E1ihjjDNijvsfU+lsFflSXuxDfKNjUiNbyx9lXzhehG7pYvcoJio93a+qMkHI
actUFaje8VtjYE6UUu/Ye/xUicBVxgVNYtK+JKe80ges31XgizAASEejiHj3R/8T
ggUM2N2xsF9iXun+VnoIFyPZ9TzI3kxlwnLEu1N4czkg7CqUrfXCmxKEjQTzOLHS
UcyVF/p7qt045yPFjSFYAxW9aBlRvaGIVAoxiNPdcoNoqA+nL0gbn6rDwNjcLPYo
YFtfi/w4emP+gOtRauoXgHPAq1AfmoXg4gHSLrjyuCBuaH+A6obEhoX2rH5Xi+zb
2Ax1oh8h9dT5yF1Ms2LM1o22pyL8tCgVfAh8j3Ij9PdqCpzTFCx8pwXTlWTIFizQ
22MtrGqPa6RnvTvFe3iflt1RbQrEFb3C60Q5NgsPZAt0C8iqGsWpDbGKjkpT8N6t
W6NhoWan1/lW8J5fGGgQU7RZb1QOd5RJxwY5lBV8+lxauf+DPn/KhzxO5AHpP+ag
4bJ45M2Urfohdf50l9NSdJ/JL7siIjCKqECMpY7fgl5d4Vt0Z2C4qMG8jURbVORs
uBRQx7GKrCx6xi8M/zwQ+s5tTkjCdxZmhlJG2OTYLIupwAFM9DRklK0uggdRGePY
2LSUrtzKt+kUXaVorE95FGbSNQ3kTdMQ1DY7XuY4ZmRDxVIqqACPAqOVocmPnI1n
W4u1O+j02lIq0DqJavCtSivl251XMaMZM1Yt2ABitTjT+5Mq8y97kFTY23PgEXq7
O3xigb/4MZ85vKFTQ/hPtk7WDu+tuhLsEkK6mc4rGSXGorUWKn4m55klPJ9OSG9G
9po6zngKcp9DtDAbOSeq2+cwTud4hdLtC1Mhz1Kqn+MlUDl4jFFbCh5xd4NBnSB6
8/0kP1noCIdAP4fknZ60qZUT6Dc9+a1AeXRbwbHn1De5DWojLzz7sYyyJz+W2EN8
LR0Rz1u1UzR4uR4MpOKMBj66GzmjGylpiGNwIRQVmsk0osHDzEHNvRdS1eHTulp9
1Se5/UMP4CJjm0Nb2ag/me0xGgX1GhQ+uCXkd3JWcLbyWktVq7X3DnHKfcmtzR2D
ZWyIb56HXTFOxMZtvBTk2m9JBkRu8wUyJTSj0goAKAZcMk7Lm6DehnOwd0JYT+tQ
+5I57Gaq5cCWCil477ncrrgbpweStbDIrtboLt447T/sncPp2q6iAb3EVFirepvU
LfIRJ52kx7f68g0GJsT/sas/CO9cs18TKZv2x9cTNxMbFfLOySkXSrgHjz9yWotn
s/kVitjryoS8VA20GT0ASV4BcIMXs77XdUwR7BHKr9+SjiIuL3InIUhntgk/LpBY
JEl8MKper1j7dfzidlIKPw1hhrQi5qY3Te/5o4K9JnBXUcS5iWL5RAVBNAsd2XUW
UjgAy5JRLs/RuQuCexLd4k4eWWG0e/VLt+JHapeyuoB2HRvdrdR2oO9AVt0tPx1O
L2eYVxR2e1DISnlYR0EF6C1t1XsIyywh+3RepAOxyF2vvLC6asIiadycnru9BJb/
s3gC4rrMW1Cx8fFyh3DIGnzBUCwrlxIPbPEWKrWNX//mRszcBM9WsbtB1kJ7y8Ss
Nwfw9MzQC5I+uz3cMmFRRa5JIUJPqRBiG8KMoxfi4UyE7+E9nCEKdsF3ca2NHvcH
JzuUIlWXl63vEezFh20BC7pjpUOfsBLLCESzYLA9V8KixpweXq8sgFBVXlVqNOS9
xPGLGtfPJba8g0yFpt1iW3u2qaQYnQyFQhCQNiXiKVS2W1Q88OC/dmfFrdr/DoKu
qEs8ykTNIXu1bRR/OsMa2ezcCmbK4XtSU3mf6Psn7rz8Y+FtpZqcfThVZdLIF8ja
5LDAdHIaO8mZQqkX2s8pR0FtZTka4U6dKvnd1YIKAu9sP5ZMiWmg+UKlPhzCodIb
KDOBJ+36+0GLShB3cz8jgzgAbXh50xRGApGqstaaA+UwsXSchZsw6x7inTO8pQ5G
6l0p+PKRVShvYi9nTFY0dhlLua+jtxs0p7SdnyJ0qSsH+XRl2FLWsk0DRGh1vr4s
xo9tvP0dicNEaydZ7gHF36pZ0X7l9MjSFm7wuuMH7/4W8YvX7NRjsMr8yivyjWz4
i6YBQZ9nckwCCjQdFCZFwzv54XS1fP9A+xdj4M8dt89n4+dNJzAVjCEodD/6zy6G
XbeRjRgMqAMMNZAENHYz1i2wupdFSBC7AX1xxQZqEQfbrDJCP6KKkA6lhke+/2WU
M/zbHyPkBbmf1qv47Yblb1Z77EFNaM8M2U8cAGtYju38Cn7YKpU09nSMHVoxE5Bm
jSgZYawjS3MAsgSD8EXTkOtRh8HmQF63tZxRULwMIGfOW2oe6ahfL2ESoVYfAOFJ
9phWLGjW+TcAM02elm5EIAAfeMtwh79irJOrEVRgNlz1uge5FufBQsiMPtpcaSvm
w1v9Gre9kiJBfqs5sCzRqFl3YpFlfUuvwsvQQM023XC96CWsynerKtQj1fG6OwLR
Q/d2ZPEFLTb1KqLZfgS3w/PdeGCvMgUH7A6k0dMMzqEiWIDU+FwObztmIJSZ8bNo
jybxoQ76JymFO/1lCfjMJtyPs8CdpfHBcQOb0t2CNJc+nqI08+vyXG000q7ncpRw
XUn4RzoSDgjoU4/Glvl+6Tffa+0l4iaMKt2R4IRLyAqoKfbDJRDgIEhnMrb7fI5r
DWENCyc8LetZtQxmUZJB7QbqR2JIkxbKp4uGQzTvUJLQlCw8NoDgdv+or9+2Rqf4
nvX6wCeEg5DwKFxEnotdVFhyqrywvvRfnshpmE05vWL40xerzBpw6FT44VXQmu1y
tZDQQ2tLWQYab7itxaCsc3smdiAECqE2CZAk4gWHqXE+mNxboSQVtIzNXSpFlhPT
oJKbT8GtelpJUqcRBoMkTzGdlT7UtnyvyNxzI0zj2KaXZAWsclQ6kiGokk+6MWU3
dEDM4CcjjB1Sz60ectccXM9rnDzl6isCMqhkRPAfsOnychXVGLGBhWmYbh+z6eTe
BuQnzx/ZOLEC/I75JqRhiTVikSMSAso0UykDVPmdg0sbjlY4LEzqbkAR1h3IeX2y
JrPUqaJvk2DLEId3jdVLmDCNzQUx2yWmX/+eCZS0iePmdRklhN61GWLiXYVdL6SW
RXtU3WLAlQWIbrvHk6z8gRTZx75X49Pt5bF/1xHfGq1iahCDnrEeNJzAx88UnTv3
e/N23PYfKbZVZAxXRJZjOCBEb8HSkDoqWo8lbOqW2WzCTjhJUyglXMSfLqnYNxto
JM+lPeP3Q1ATR1qIDPd6VPnhTD4KSPha74K3vLMy7seevHbn9PLQ2IiuORiWIqWp
D95727/TVFymsR9GYazyeqvC5TuQKvmC4gi1uh6zlSUnOtSREwXCNgR4gOTCV+Yc
7pZtz4oceiyzE2eT6SkCTwiRtdbA+vxBe9yl97oPrOaByl98JopIEAiwzOn6trzy
xXBmNPGbgOZoinJ54Xg2p6yRMQVEPMsKm3shsoeqkzbgyYilpX0/bRjHLfzrUDmc
hZ1VOilrYfujtXNsyJPVvk1ArNrFeqp4dkxwZBYzTf0sgHB0xt8Uco3TtfN6YLk8
j8A+CpVC2r9NNObI7w2MTxMjJU/Lryx5GsqVM6iUA1r/LYZGASWjQik+m+lbLs6Y
q39/MccDS+u7takt2JuxCTfLdOxfesrqs8Fzu3zvFX+tXea2Q68CCgWc8LAJ2943
NRhDmb+jIVB9m54jgOK/fIPYePFSt2QH/s5FubzQMmR6k3FUGbQ6tSQ+tHoEhJH5
Z0wqXSO8mUuUiVU9HijcUEDGZ4/WLFAkmJQOKi3WCGkoZrYF+/EnYt4fPRhydNnL
MV1nqkE+uKPHumXJ8TEY6+LCA+i5TsdpILpg1o97BB+SYD0SQ7iCqBFrNhcwnfGQ
ZPjO3HJAvCNer2v5CwAoArqqXjoPSHdr0/TRnh9YDyUoQ3TEE1B/ikbacRb4CiBB
l5R1KstJZeuG/dQJ+roYY9XbLYfAE8DazX53Df5XfPlG4QQs8S9RqQD2LzdZmJrX
D7rThgMiIvBb7aFgAgp4GPkvgerJiFykwlH6jiKW/ibdQ/HmJpQdGNCFlVPOJ5Yq
U5scPf6WtFGScq2ggKL8l8swAiuXMUOaHvY6uYa2IveMbZ+VLMDF0DI16eHS5YJU
XU50Sb3gGvgvqo4ON9EUWhbRIfmcwnEuNUOJrfHRtsE5dWRjm/CG9WSPBql8foX3
5Ki5XI8RPProtiQRF3gG9wNjKOvquRVJHy6KqkrGyCIS+EY0XD8wdVKCSz0Rj1uS
EFnSyCoELAFyjalPu3MTnLQKFoCikjrAFUVS6fRalX7DYPASp5xLHIPXdaSESLUU
g3p9dRtGLTB6bXIMq/NqUr+tfUcGYN+57rmIGi3HPj3ayMwoVZa7TEd0EoVivJDw
ubs2Fk04ypChGna/2KFYZ3n47BE8uUAKCnxMG/PP+IYHIlPQYBcEA9WNSzvt4cbf
XDW1M4lCenNJn+QvfZxdl2qqOZuZzB4WrlduaGgYoNE3bkAup3Yss1z4pTeh6nZS
mipZnVvlqDW/imbyy2OKXd3pLh57vuouDDGP62e6KZNjigIUOBRWiegGGZZBj3NA
MT6HlHCPmux9ykkyFKMyWiFr3w4L32XK/nX0b9Rupk0pjQpXbnmU9s4tyQ6b94XG
0hPuSkoe6xb3RhbhCaxo7dU3FUeiQfMAGg9crmlMkEeBA+TMvkUeVOVqH2P+95zt
aZp96zsgxARGEmUY4SOn0UER9RJF+xcojl/d+oDt+LhoEbrHHm191NJ38gv6xROd
XfqlniPUfSPGC+Lyw+P8I35VyrYHIGhv7xWZi0E/jJLA125LpC9ow0NHR0uxLD1Q
XRmujKa/y5Kex+g1OkY6godKvXdoWWINHJAVjc/ihrbkAuxeEzdeI3lU1ia+yVUV
d72bsJUCFJoUGRG8u8SGtPDW2uTUPjU5FB4Du9g8lvL0LHv8A49sOo427pM80xnI
mReDmgVR43vbBXBh3Xz5Y0H1RMEiOByP+ilzl3eYCt7bjcfrPJsg0GiaYdfuVbxk
Lx/JLDAldfOi0b6QSkDXKfAqiTKjQGRRy63CSpi8HNtpNUqUNHkvESZi+vkx5mZO
59CuI56ZTCFTkV7GvrTeSqB59juqkv3C5gsIQMxbf3VVXZ/NX3I05mWRXu96px1b
q5tjNPMAO6BiB2/HZMgnw8/IIvctgu5vzLpd5p3nA6ySskf+5oAy8DL7+rwlpfMv
/lb5oSI9iGKPt/gtmM69pWylrKN3Ype6+AGV5mSje1NimkVDCmAJjD8D9JOykbpl
EieFzNU8GWkakWOzlXmFOLFqVedBzr++OeDEmF8hKXFTcm7Fh1m5Czr8DVzzokdD
vudhPE9I+fxsOatPWR7I7/kvBy7ZihpWNLnjZ1N35du9mIgbYqhrZPbUwhK/Nckf
elkWCUJK1xHEa+omdonTlGm2J1sz5pYpprnZEjV3Lfbshe9N244tIzRxTUeMnyi/
bGZSyNHcsH401jEF/Oa5B2GBBkV4hUsdTbqoN13VTw/+iqw7z319jqXT0A0z58AI
r1YK75xmezJT/TdkDLgjI0O2HwfyQqRQ2MoNRX8nCUj7UGYU8iMmQp45MyUH8Mh8
H3YxLkV8lj0IhIRTrLg9W9LkFOdcorn80zTcpI8WMopx83ypgh+0M0lfANv5eWm8
ZgxWOgxCV0GOajkP5wDA7TSMm4UJoZEYk4y4ikDZgFNTv7L6QKWN/o1wAcSeFuiL
OAF6jQN1E9wzP7Vl349dI1Vc7o/hNYhQQ7xynP2BTWjvZL1JuXVUQs4MGBqp1sMi
Uo3Kv5tv6VTo2qmbIp4J+DM7S2zKGrOP5Igg42vtufyTgbuvKxsRszat/6OfCMtD
2cuvc8GFV1BwgUO+KSE95k4HQuOVUsq8KRrgPj8zzLSwO58wUT78tYVunVIRz8tc
VPst6dgaEvixpxVqrmLwQjGbws9iJ6x63zrZwCqOYYyBeheJfIqkWAO++rnVkU9Q
jFe3mh+mhYiUDHsnAvZ5/rGyEC2+CcLGpoqdJJRTH+nyGZJYhWEqWobir5tbL5Ow
mIHtzYZ6Kjvl/b+SM5ZhdngewYoRQ+qXi/6waygUizF+A9j9nSQ+xlmkZV3RNnni
CRfXGcAJ96xXizT10B+I7xaqj+nzfDPV/B12WqUeyiThvRG/AHDQKSFi+5pqtV6O
2Ip0I/v5LP+Imqn0NcOivtWCYbIl689zK+n4wJYV4dDW72EVjU4rSfMnVGwdyWRc
eCYrNKKj+H4HasKzOztKDyynzCGeC4m4Kua2J2Bqs07gxNdRbpU44jQIdunejoPQ
sexIB/GyR1uYE/G4QQHUpM3/6XCm2EQluRDZc2m3o63CssuNreDzdzFB3NQbns++
5vHxHpE143DI430AboPV2dLP3vlQtiznRfV/9SPvVp433gpycQKwM48tp8O5AkU3
/QojHy7k+IfWf4sgTAplqzyGIYPtGvHzYe/YnhgcRuaglid6NKfL8oQozTFKoTpD
6iT3osZ7D01SpEyxBLIN3GarDukMcXNmo3dxkOisLnT8pGVmWmzm6vxkwMtUUfWI
O+Mdh3e+MCEGtDI6DHdNR1Vy3AjZYod3Z/5Qg/jmf0M5zrgVcW9ujapyTZr7nP2p
NH/Rd3h7xiPjq6fn0YaFXeI0rYI5Bf2nBkq2g8LsQOAC5Hs449upmuNmD13gGbQb
VU9spv7eFN3sZNNbSJtqXqkcPhQtCPNmFoK5b6tmt14GpP5nvQdwMa0nMVXFxhv0
Zwu6NSMHhRF+EvBu7Eg1oOzRxvUDvqzhvp12rSDBhtvAAiv7lmIKS6cL0IjibNhG
qg5nU2eMQym5YRgwuajHg9EM78GGyxLqyOSBAnLOJtpMEnA+vJzzwPh2rAmGKzpl
jPXVrS8ilQK5mU0jpCl/FFCKn9/bk5FhAg3evN8i6wz3uVhXxMUCCQcBtHsFApz5
uKjV12m0AW4nMdV1r9ugtfK1rJasRKnILt9rqzvtiPfAvBq7C6Q7YNp7x7pR3MQm
l0HHcvUnkVwRhE6WQRNdkrEHbvTYJQP2pSpaA3YQ/kTgiCWuwm4BnDIWFUx3oqSL
oXd4Yc2hJnhSLH7hXAsiPWhQlzzacKMzbFCJOOLKQ2rFg+l9FqnqmFRx8HpAOyYd
5ANNCtLz2hFE2MKxpVi1+vCslKqercEdEL2Z4pCmkW8E59BbFYHsmtuWHbLnFaAY
mQ7COAolzplypJzsKww+/PZg1p99pvJrvkugUoJr3MP9RUoMT1CJQqVQE2BkIPgh
CJfVaw655cFHcRMR5pNTJ7TSBKn/HJDd434L+WKFwzIP8UOGWilRiGHLKtAX4Ms4
RIwFOiO7FQkLwE/7ElgaEOqIfvhdYhLrzX5Cuh4ObHChXfqdFdn2+wPFawfwdNY6
D3ekNmWaxmlgWepualSF+LVhSgzZC3xn1fXZ9yJvJHleDQHmm3DYM6zRPWtNn580
whc+NurOQPLyqLu9os23naMiGKL7Kr9YhHuwyLNOZo+CBUMVYeoWx1+ireik8Os/
wPMLJx0SJ60s+n6LalQlrgZUPkQ1ylaa2O4djnPF0Yd+2v+cN4KgpXTvyiOe9IeT
0xp1toC1E30QgoJNZnXCegZYpkEVrhVHDPA06LiSnZ5w68kPgiqEjQOdeQgTKqWL
0mmsLZn41drUZJBaFYJPh95NWbEU1Uk240X+DFsAHSyA1jdPD6H2Ac6A05X+u1Si
5zSfOigFvOGSyzrbcPI/HquhQK6pd35rYwb/kZRC1u5RuxSl5mcDhEBS+Q8Hv8E8
LRQr5c0+txjrlGLsUk6sMbLwmWHhbB8kLasrDa9l/+N07DgM5E4JC386OnIY/SfY
6N6q/Jo+/An28cVixEn6w5EG7DSu6+R3Fr0gU1jQRblfCjRbL1PQWySxziybBCUh
uNMeQsKcBwYC9UjRBX99vMGn72FoW9Vhhg+4Wn1y6wkYuWiQ4/g+kLJy5aa8bZis
0wDFboa5uma8HWtkT+2d4OturrXMzLggwn3jQnNMJzzipt3likumqM5fpRy/ourp
rQXsp838UhECqEl563AYw6D0ayQd5YI+YfTjrp0bMNrZVG11QXhvDQn3k++hYrmM
5H7sTT79L/RfnLbONOK8dnKMCEg9fMn+LIxXBd/s9f9IGH+9cobjAmCCUNhpS+No
Any4dZ89ndpgmMkX7JjWvKCuuVFGLKZL480KtIt22x08YT1HH3hVMsCHOxfMKNi8
HCCqvXI2x/ESOhsqRPvvxcTEiobqJ56QzHhae86O0Wn362yq890DrSuWzRMcmW/9
IRo9d6YSqofGrLkSmyVPgzdMOEvOQaq0JTukrcQxrVG+EeiPDSJ/iCbmBGCYe1U0
iYalw57PVHof0skKe7MKH3Z5yJVSmmtZmbYLqsIUFI1YqyVjJK+XgzY/qWBPoAiG
UPG0utp67v3K7ZB80ya3Amck8HFqKCLRHJ/YwjkNmFVMgwottIYXm11t9ABZ9e+f
Hn4QnOqM1N/U2/2/Hv6p3XPLYIgjkF7IHX7NYxdTqYMgk7JizsnoGdzrIlwPDSvk
LDU65RWHEalUi5IUCVf4zjWOob7Fm9XEgq2jGYoDNP9r3aajBZpzUKzWBooT9nev
fnD0UYcfHoyrEiGq4DIn4kkB1a1TdF+6ec54L6U7dBdhePGuOeL8mzQnI5yYdzm2
A2UciyF/tVxdDNcwa9Jm2pXuLwtsJx3T+8IaZ4erKQpnCWWHmU6kZMQa5hk8dLuh
erjKxR4tLTM1VIUhk6Q85RFdOxYLNz0pgFAwXO0rY6ZjuoCZP1aLwIfu40c6xKuO
URnDIO3uEN/hLph48SXUfy8RLZsiKzmekx5lzevED4sQYyMvgGS2mwQ0rSli932P
pgxoHGvieMeAjxD2aPKD5GOVdRnIP496l2yGIn1rU32BRSOTtDJ8BqKEDxk1/5fl
+NMxot1wCSk/M+HdoBkedMz0ltnZbJdiBUm76Go70gVEp51Yuzy/ikLVglAmSkW5
JvLnNxDrzID1+Y8EfebT70P48qPjm5bpm+3u/KUZ2jIcIZGq9LJFlbWGriMePs1+
2zmoeeTSPQFxHknS864uKoWOagu9gSM4MrRUf74+1m0KrjfdXTLIEL0DiddvznXd
Z6Il0eqayirjzOr8w35Wbi89Se3tApJcobcFcZhyi9qp9fmH0aVRNOMLur2o06V8
cbyM03lAhdmOG1EqzDguoBwh6MslOmfQ6NZnQo9ShhyxadwAX0v1eG3eE6a2bJfw
YttaiU4dRUiKRVxKr/rc7Cj2gYFo4bPhI5D4DkwhUaTL2Im0gFFOPIv+oHsfxYgF
Vpdxc3Rs188cx73QUFjJaXgy5u2GgC2t3aMRzeINUwoaA5UY+/L3u9Koq1NVMNZ9
vK1fnNGYWvMAcR+fDgTvDnwFkJ5Z5hJuxScZ/rUBbpmXzQLzezPiorqyXHlabLNd
kNC3xl4z6VqhxkTSxomeKqQd2FvnsmNv1hspN8M77eUZzofZjo5hxS8ACwYnRjIC
6GFGUCcggHGJnRJPasGQHCu4mj5oPxWh2AX1EtyDdIPRcBCIb+QR6U3L3kNiE+1r
p4Vddqi96TJvORKUQqU9SYoXw16d3vL1sWyzdHYoPXSDVQm1PTjJEYzvEGHYS11V
tJDFQLSUcL9yYMx+YojYXAvTx3/EbyhNgdZ4xc4Fg0GrNU0c0boIEITypirqy0tt
hcLwp476ypl/x0zJlikDY0JsAduYEHK5NzooIDYeje4GdwPF5iFz+WgAdumyPZ2A
MkXXgsnr+3Q3hdFHWRSGJrtJ8LtI0P46UTbp1MNL2V44T1bWVZ5cNrj/NywPox09
6pedC4w3UF7mKLc1ukoVVSUkkNzzElpNsJPBCZktLi7tUlJ3hNKBwtRWCg+t6s9a
foXcrSUrfTRF0+PNLKO5/KfjmkqX/c8fdMCQwGRS2dGrJAM//ZT8CYSAAoqKbvN+
MnbBXZTZcmtngy8Xpo9qjCadycrk3GJQ6aJ8Hl0sXtsdF4jRRwRE51thjr9bKYpJ
5+f5cvcRcitiGH3sarBfU1H1CPcZchDDKcIZ24g9/OovVVb7wQpZqL5rQ+cGbduW
j+2LXMsp6pN3w1olFVJy/DzTx3bW/OBdWqyx28Jn5vTeiGGWVkirYQc9881+g43m
g9KoBY5OaRZf8S39WuKVDokqHr1x2m4UfsVJJ34LScpCTqv6MdfuB6MCf4BE9z4Y
9WwHK+b1kl4qq9vB1v7cS7n0yAuRgKLbQVcWKkk+Fj9NFWqHKpW79H+6KGYFYYUH
TITpFD01j+LNPKVdRAK5IdTuzC4iZVcNIRBnYn5TE9MGovHo5NPZ2Hnn0itbTFEl
+wYjQ2v1329Jyc0m6Oy/yWUe7Ipe1ttvpqqsOBjOU19lGl4ztiu57kukHSfxkSh3
EgmP2tJIebYgf2jkn+sFqWRZmLcm6S2/VqBF0YhNRg23WrW5tsPbJdeZRMbVoOcj
1++QZfMSBZT35rUZhrCmjYcVCbAZ1ZEX05sN2bhvHVEcMVL2Pfob/yfqVlddUsXl
XHxlTcuqVpK0A2E5h/2mV+AHYdzr56brhIttt8NxaEheuUOqLMOLiOJATBtrrLwJ
SyBcIFgafsKOthYXKLZasNR00+r2TvXLpaJnKdUUvvghvZRKGuCpwNJST5WDgCK8
E22Nzifac35MHqAQndcBkNhBEHF2F6y6EkYu7P3qZym6twHPvKml4i0A4zla7XAw
6D+QOrOjC3njdzndZaAcHo7bUUdIIB2lDFzYx1VdqLHIA+Zqt+SFAeKjwLJwvTFQ
M2SNnG7OBzRu0hyyPoOc8VKq5fKb8/9seAYlHBHZWdDCsL8NJJpMN/TUDdWELiQ3
zguIJBVvlBHuh82KPFLgj0ysMxPvlqB2r8KzSxCRImfuvtPAApLQEchwKmEab72q
P4yZIvOlEFbwyqmtwHeXNIAoTtfL1pYZtOUeGomRcXPhMn1NhhT70FsVZ7jwew5E
H0U+e8ksd5qP9cSFaQmdPtxSRopB7wj9vvta0npEV1O6ORxGiMP5LuqTXMISl8d9
Myt3zUhJr7D8o24m0nYRpYZlRdM1+4mhPOi6p0yOpNn6bU2SJ8iucuZdVWYwFI5y
XD/Jb7UndzuuBCxShJkkm1qo3Ll+z5VcNsBHas5A1rH+P/uEAvc7Xun2z4COPgyR
/qUr0ZGifDHWqClQpXg88CM+ert1nqfEKwoSdpBTVcAs0mW05+WfIUB/92wyGM2J
QASriSgOckiW4ghR5tg4bCeL+TzezOazI5picYrFH7+XrUXSx8XZs8eoJzxSKjKB
nX4KRKDPjk9VL2lnvvxufaQ/Sd/RVvLU41QuUQPSJWfRMgabYUwVnWgQ8X9qLhca
MoT4SuOq2tK/VINZT+HN6gI2TKZpmCJGbfzahDGdFGG9qnysIvH42aaRl9RdglAJ
USnejQcwOJyACXDyzQOUGutIv5qrL5p5UD1piQz7v+/W9U6QIvpWa/fGVb2Y4kMq
e6ZzpyBrgmW+OtYT9RXPzORatoSP9PbwFZYWNXtaZAY/n2RqUy7A1HK8irhL7Esr
h5NVp4IaVPxkKPrdof+eDPUSco5eAxtvh0Cb7/i2LQyQrGimrx+dibcKORmvQF+V
ucF07UwszkClhJypMMgkrOFVbclv8ER/+mbGcvJqO9b/I+kSHg0D8JgODtMh54VT
eCW6pRsyq+dGpy1diZh8rlw399wkZWR/s6Nk5D851IbfssqEviVgJOwxVnH7ZniS
bnA3EYyWDFyvFs7ac6ckBxwCoC6qhbPxAr29ntWPCjqFgTDlP2RRfs13vW9uNyRo
WasRWPy+Xft7Kp/hNey/9FiO7WQoW9gHEKXLpB5Bzd8lVNheJ77cxOHWzGJaPrt1
XyFU63/eqtnsM7/t5hl74sgsWdzDll9HyzpQ8J5qx+Kdn27ZHkHtfEbH5vaC39cJ
0aEe21gQI8W3dPn+SlEUX8wBYGAlAHmC784pcusamhP5taJhvYMkegGq7Q2Wz6R8
imOi9pxyYrTce+ehRO2dC0xfdl6jfC3K+nnfe8GtfhsnquOB49om3m59DyUU41BP
uzeeGz7noH4hgbjD0/6SlMu+hlm4QWIFAMezPYNAY7mWW12s79XzFmCOVJR3FdwE
dYzFSMbhvTdr143VA1KqXNqOvwQ2M4UnARlxdmfO3+KV5kOayTibGO5ZS7e0Z2y0
gV1MKL9NnEBbxVerFKEcsIH+LGeC4IdZfxb0VASuBP6wCbQ/fx4FPabM5VUjGY6n
CTTvySCmark57CZT4W8lSChoNKdlFOC2x25NGImPKs7cDWqUs7/8kizAn8jMN6Db
uZZflETlAgpE85xo2aJasUELMLERudjG4CjTIL6WgkZn8CG3DZrMo7tZ9KRf2Tdo
GZmXr3raJxcPQpL3iRK3UlgLGwip2gcuNDQA0CaipfSiQpo2AJZgBB21lcoGmS+G
vG5o8zkRY57Anh8TaaFEhxbcuRsq1YeGCa5XGTtrtzpnuc4RlkcT9R/TdPbz5PO8
NJVSlBDjq3AkE+g1aYlaemnpK3KF0fIF49ZunD2w59MXeTRgxF9GZwC9yWj0ZKfa
47xaRvkgNGparm8NS6B2KJgNKMCRiASUVd1sjdMa2u/p/rRuIl4j/vASo1pwINsl
hgXXGw4+oiQefD2tvpD7OaBdwYfTi0UysaPzWdLCUYOHp9tjHmuWODoMqcdpYvTW
CUatHM7XPTiyuFBDzUZFJ19tHx1t2E5y5Ibzfd4spIuOBAPZmnaXCZBa0qpPEAOB
bW4bniPQPv1ZICI7A9Mlvl8/ytuRJpoqWteUsNhUY1Cvdo0Yv93/+ipRrT/C+/er
+LsvI7jrZy1wZyeDJlOwwTnsX0GRkPC7Kwk11k+fwoVS4aGTzi2hJCLNFR7zXiH4
/Sv3DmfETl1bBSr7CF/+0HCg3wcqCiy3QLlwNA8f9Pld+pye4VzyFMzFg3vGKSCI
yeugDVSdMasdVGd5jqRfixlMjoUz9pNuZ9PD++q8eMFRY8iPobdRVzfvdDPI1ggP
btiAG5SENuoIAfHXb745koJzPS6lIXhBs6YXa7ttX/Q7F6B2NBcvBvtDd86khaQ3
WEQ2u/j8XN3hH1MUskPc2jxerrwf1JTM5fa5u6+ECxEirNj/Aw62Tg3hezudKKHE
LTxm2ACuuGUiSd52CC54W0enQ70TdgR6WrtVCHEK7949qeDhbsBL6BHDkIyiZvVP
gGmsR4kB05cLPJQx/T5iUuIV1Afgof35LOKMAvbZhS48On4kjNSilP4yCXI8U/iI
UY0q2wJMkyBIdHwrirtNZxZS5JEvKBgBOiz1yI/wKrQxU56MMTppePl238hiigaA
i1ThWnjcvm3THIew//e8H0aRRmgEAw5a4ZrGrTEh+suQe152XK0oT1+wtmfmmxHO
WDJHpV2EJi6ciIhZqX5Z/ypVV3ywf4C4LwZSGUkxAv8PRafjUJ0TDVG8W9p9ghgj
ss1s3K4fURpXDaM1RSlQZyW4m+Yg4V2NZB4uA9wIMKMqN0FU98mOqMd5MZEeacEN
LLFhQ7/5Hk/9dRK/yv7gLMs9zSK/KdkoV5eD5zaHWwxrtsJ5dqroukIW5doshXSB
03gCfN537PG3T8R5nnriKAEBxdKxlMXqwnRKue8qDnbHvrolSuXkwjlIp6XO+WWI
pqOyFS3yH+gG08aPSyxIRCD8Hdxo5niLHTVcMUGeolXep5WOXqhjIvKp3fvo8flM
unfWZd1ORkSvEXBgxlmqGIBZzF/LLZOmRgLrYcdJUDfeelROSOeDRk4a27NayKDh
bZK/cCohB1TS2NNiExHCPRqpIUYnq/vNqjFtuFgkhp5w6t9BXMFX/mpo5dMWcWWZ
VVw1RPWLc7YBKq2NE6Vd/bNQ333GVk6OCX78XdEqiyMlLarU1ooH3q4MYloP4p7z
wEvYYN8UR5Nzlq1z9d/YXghmQ5f52HB6ZTkuhjbzMcTm6BGgiQZB9t28qUCiSqJS
Ge4GVEYZ8BbThmEFgN+izbrliqFjoPOuoK1dLLAhplUNLVYi+0bKfLC25QEMN6wc
5ozhtjRvErswsvE/nDwCr8F46V3ufWK5Ey/Hu/yPF2IQyCbi+P2bJ5/NW/c0nIau
n6MDpq1bOZkOL+kIAoyVMqFklZC4W9TENZdZ1vcuafX4W2fHTFU/f1bPCkUNS76W
ImaCIO7ThMDfGYoEs9lFF3624U6xbvcPqldmVQXo5/HfRGIS14yfztybR7gXtF0E
5Zc9xvgKGR3EDZva+BfUHh4piFYbvxT7cAxKo5ycAScKrE+eRtU81+OMl/P3tY6r
NEOb+1KJayhM1CLzHfJM38RDJJ/IbYNYigg3FC7lQe6jyP9+822uEgsywbGnaSbL
coNNUVIURuJOe6weCgiuGtiL9KzqIjGpYRqZpTEGYlo7fTOtl+lniPHjTNC8J4a8
i1H9x0FUXD82JY04Q0myu9KxfGr1+xFKqshVrKU37rHhHzZymVxr73f83BK/xtfP
PNTuXuBm92YwsUnqV7gb1sgXRtcKYCX9du4yjBOpx6ej7ZW6CGNz/42f/AYqcqrT
4RhkYUsYV3/nT8/PsLCmPOaYSl2/MRMJ+c+wQ1jJoaxQ8El+5dzBdAKRMiqEqmBk
LVOBN8/O2x63r5oOs8nR03yH2YYLQGgCiaDKA8ReBB35bamKwOuVAd9tuilRN5EZ
jHC+uu8TClfWxLJbXOKsHTkedhVr4knlxLkNzP1UTevPRiKIh0tmBXED+wuoT9R8
HbchRrfrWLLxN0bCEkm8QK3+Pd3vexqd/1HwtlkY+pQCzDDMdDNl1V0cto6cHPaA
ErYAGfDugp65S2qEFC5jjSqrBNsEiX59vX0j9xl7dpnrfJtiVwvDvUpzyoiDOX/x
CcPLJAh2Vn5j3OpMbHBo2tkizEYAKUzEwEkCY5/XT6nfq6t6Iv6Xy6bi+TMe6EJC
wG3ZjaNmdRbpC4qR1pzlEgr87fu7Z46paLOHOdn3gqz2lDiTxi1fwCLfEY+hS/iz
bf0HY9sXu3l7RCxUgkeYvGSN73TCu9nswOzy4dBDAb3tsPASGU09jKu0bm0dYEiv
TpBcFvzcuW/odos4dyu5QZp1FQRMEIv3fIdb8332lsdFO9NN+p0ngVRG+TbDGjah
1gIbZcDKIpl4xC+tBCiiJ3SWO+YGBrbgqMVtutfBmTDR3QI4OXdBSuAaJTlmgYxh
9+6eSV8CBon6gZj4VfhgDg2bQkKqxLKL8872gwHPtoLZMfCHdhfzQYkLibfL8o5W
4/D0vahy7ORQOGpGVSCw3rVOKyuu/h7vX8vFfwEeuKtQX7TbeelBRar1sT5SGhxo
bPRc+5SfymifqI7Kx7bJwmZysmW4ixsLP085ER4U/BuO6MapfMiInkvBpMWOniu6
SZ5tlRUmFE7KrGash6IdSsOhWWBC3K+BHRIPI8U23Sx1f1XeFO8F6zdtnA8JvVcJ
fh5vmqrkznV8n98k7YLcTxFy3kPlpYVD+D76eOdPsO9T6iBVYmTX5/I13cDgNncu
uonMBT6JsX1wsge+yEhiXxp7MpdusbOsmfntIxEHHQFg/gkiCTQZq9lssa5ZJHPY
CBN283P5qsNaA6JiBsRFpNjlBGSVws6agxfnGBaWtdgKQmYlgU7/MDNp2xllxQNq
fzGL89/1iUo7drXEpiAHB2HVRhr1wTRBXVJ+HajgWMME0Qig9O3RlO5JipTxuf8q
U1Qz3pVKwdJfzV5MzofjTRwoophTUDILID/CVVLkbsBB6PBnGrcEXINt5pIvhCCL
+rJ1M/Y260SWqisnCL0G7M/Y9d4mM8+sYUPEGgQ+VCO97P1+zBMxGQjxbcZGb/eH
p8HBltHUtwJrRAlgcpyCKcGQXzWIY0bbnIiR951h7cPuI99G/kSDZW8vlDKkEkD6
M+pC9xrFdXpTvrijMcGVX7SoK+jL3YetbQPCReBVPfmGlaqlv53p/l6gtj5NCEk3
4X1swpYqVfxV87NhlMa/xQtPeaTSd+znK4Q9my5weH9VlQIw/unEp6GDhqCTXXux
mqvucVYUFyHMebbLi+N4qYhO6bBycPgTAASREeoc6P0AhsUj/ipTgkJd9Hhytbi7
spQmCLsW1xFEoJKoB/O1An9ZdBtGZ14DFmt6fVp6RkX/5tidDtCuOwo3jgrZF7P1
tjSUSwLXqGFX7++STaKWlCLU2RDLUNhmsavPt5GdgAeov2WD0bnJH22BuUqjDo/b
PSatVYFJAxkPkDDs/ZvAanl/bTOzPTqllGz0duYrQqyHJOui69oT5Sv3G37Z69m5
DP2op7YJ7hBGoYXguzUDzMB3ztcT3C+4skRB21LPcwF+DBEvPmIa2o3Bpqb9HoK5
NRhKDoSTFqoWjqpYRL7XKsh2qRIyMMeQEqXPpqtRF7lO24RKc1aQ9Z2lJSJriBkB
jert9s3UHVSYLyVC5efvkMKIUx1ESfVVUA2O3wl1wz0600vDH3IhY6J77yEFzo6I
T/zSygOV9Ss+w4Yy11u6Xai9rek52dG/SZVdEip9hHr/HF0+xLlCwiaHUOmDzAOk
hbhbdZ7q3wBepx10eNmvafxQu7LfHEDzDQLBjibErEZjkLJkOWMV1dcW7A2uK8YQ
Va1XvFemSoWmzBisXrcC+qIOBlZbUnDzwMUt7iwakKl1eDbBogxRVk2Z2SShGIbx
iXSnThzgesPx0DifGTUbelvv7cPBtsinJFMK0bMEK2D5xyfvXQxnJA+o3HYhATwn
tmhhukppmh3SlcXRw/NlqhFbzO3B/I8wtl/II1Rb3p6DCMcTxY9hSIRKlZqKHI78
m4zvjYT6IP84226DDxIRYEBx90gFgxMKd2DfF7RG+MDO9YeFWGljO7JAV7GQzdAf
BUN5H8wxyRSW9levNmraeYAlePCxy/7AxDQF60RpaKh11XF5Du910orWAE1Rzu3o
P+GZm/sypNhUzwvB9K5oueYtZKELe4s5tsI3FFjFsDF7zqlANJU4ClziexC9Vc+T
cthwgARtDF+l/VIYASj3pneXzp4AMsQZ+6X5Q7EVPa3U9xXN22oT4cciy2B/u9Fi
yXQflry1tjeLbU0l7JktMbEkmZj0oly7VYwCFF+Y6GjVoLTCdyb9k735hEnsggx1
635djFAGvXsIim44oLznMMi6TfUpf2umV9UFF3y5qqLHyLst2mx+tgSIo1Qi+nlK
wBsHPDBwmlUDPwdf/Pb4LTc9RJCcppl3OmG97wocHJO82wJSbBY+bBLB3DWfYzW7
dG+QkceqN/sj6EJbBu9rseDE7rTfst9ZODwC0MQXJTRW5lRs10F7h4eAK28sFK37
6vFNg1kOGKOhaNrzu0SloxvY57O59W/3et4PzKs5RAkCYDCuehck7SGoNtoU1+Eo
Bi+yNNKKry5R4Vzn9nN4IQnFB/C8R5feiAydCS1VXh/rYifth75h+xMmpiQTsrVT
wj5+CXy3h1OtlwUpsoO2hvqSpW+12dxTT8wAgizc/aiS0OPg6BJM3eOAvpk0XwUX
Qou9THEmemDGkjqV/vMGbqLXkQJd+Ux16vBYxTefh63ubA1ZKxwWfwoi8xqfBrrS
ETHOK2TPUnmX8H5u99qKkZvUcC4Fl+KYkqUCkU72a9+ZITWEZNh6OoRguOpO+H7r
pi2G6q0FsBVwtQkRYePFZXLf8AlgXL0PwQS8uAnFkpnhURzAIz8qR7chWKmtLQSO
bLpY+foODMNSKwNbfbfEJy/iYQSEeE+iWtZypPTA6Ylw9wiykl4OXZlZbQlOyRU6
EflM8JuK9A2RyGgnWpXMRaqAOPudp2uZ/H5iLmhpNSDOoWAJlDRQWWGKn4LlHQ34
ThWdRPJpO8YSsOm+qdMXaNQ24KgwzecxkdEszPT7gE6ipnG0rAlt1Sunx4MC66Pb
XxUnWYiAOLI4DQzWP4ehPhxWYG786owunwchYD19h6uNqBEOArHzpe8mumkvz0Jr
49fq9drMBGLXselrnOovEdy+oLbrBBoG4CdbrLKqrk6POFMHGXaUcoTr32iyYEVZ
VyB+jw7wqN4bb4yE+rc+DxzDb/LnJdLSsDXcwRiTuHx6/OV0qlXLBD4uSVwrPOTZ
416aNp8/PhapvPEF4GVKp1+Bx6Wo8Mmbp+K9VXij2uUMS/aLPsx0gqilD2Y+fNje
7Wyxd9qogtFcoUxkMrREcxJCyOcWTVeLm7INDPTFVtw8YwT9vd8Kv2PTDfVwrDfQ
s3ygN5GPfynWsWD+mdPwvGC7gHz+gwLl2Qx50tZZvUUmgXZtGfiBeQduIWrYh2Jo
mTrtNNlPOhadEQezGsZVldol+sDghi3UQe7jgBF080MPmHUVT4Y1LZjOqGacFHWx
Nvj1Z/r0yCQC1ANg8ABjVMt+ACfC5yI4qAaZsoI/lEQjIUsDIJEuBvvlJgh8TAJM
p20whHlK86bQ8g9dPVuNKjPKsmIm5H6XRdm+cHKo9JawQytrqA3Ghdrg6/Q+4Xb5
v1GmQyRJNR1AaqUf9afCONtRJK/0iemvFpVEqhhX9JM8vmpQTKbjtWWYc5ME67rB
ERiyQN4I7aDHdmGou7kbbw+XvxOo2vh2sjPcjfwKdYRZTWOSkO2coP+iYYj00C9w
n5F3I4mF6sk7D770LyRYqYXX2X2XBCBqUPggsT/R28jCYoIp5DiymbSLruIR5U0e
zxwBKbYoP51efohVr8maJHMMz1ZV9kktc/nO+8ZauV5nFVpyNybp+Fij4lg/EZIs
Y53GL2TcoT1+RLIH+1s//93x12AoEVXvrN5jMImUGzGtlrVOOo85ftf5yfhmlqmx
7wjI0FFZOUARo+d+W2eUAxujOLQ/nnXHA/oMWTA5Zm8uaHU3DsdjPb4OnChHKBhz
relIf7sZNbGuAXUBqHbdM6hKJzPV8jzHBvMt8tmEJBREC4FoU8S73cGPp7m97fdX
8dlDXl8acKf2vxB26R163mNiWDViL8DQV4ldo+M0bsx2s9uQww09IbCoqhAcvnd4
AhuY4sz9OX0NhA7LY2oDbojfjOoacmJuZ2sZAilwb7aMK6vov/xT2DRP7SnO1L5i
D1Vb2OeAcPhQoJTh10F4N4Z9HFyq/g0ZUqRRFDY+f5Iwi1BBlF+U0pjmeFePpHVm
l1eWeJpA7+hXHyIo8kT0i2y18+0D6hPSZdDuiXjkmV6h51CS1hQIuaQM9qgiRxCG
ESJ6YRFZ0WO2ogW+oyPtKQU7aX/dpL6GQaSGdwsm0jXyelvse5xnuNrRpHG1que8
lRf8KwBLWWbAbGXnA56F9Oyb3zDu7RZzJ+ht2X5q3PvO060VDmz6RSYBNQJhUiT2
1dxnc/XHYEbFgkny153ZZzqjkt0LNDM/LNkSEL8WQWa+c57N1PN7PTHwaie2kMsC
DTA9R57oUJGRChAf8U00qbZHPeFOLiVFuGuxXrO022NTmqfx68PjaB91kNKocEue
GrKEqdKF2335uHdvoS6uZwKx/NxbchHMOSYxJhGlSqTPj+kFlMgtkXsTg+Q3Wz+V
dMj6Wq52OasGyVVktK+hWLtZJoX8/r+m8oOkXzRrQtmXA6MVhB4Vmtn2Iel2nBzm
VPd/kfK87Bk4DQNbHYK1lx+3tV2gWlTc1Y6UDolmXbQKyvUOV16edCSfhM1ChEUq
Hk6br4cMjICN6hR5S+Ds8G8YnCK7/tDTvvw+fD4aByEID73tggGspFxebRMiOQDL
lDGsnMynZnu1GfRxEF7/0VsDpxgX6WmXaPD7nzWCLKxLL6LV/BaibqC6t8Runhdc
2RtGanBDgRT6BieMPjyC9Q74YZsPWFQRkFQhZ+erv5dZcKI2gNV1oxObSdtJi8XW
PAb2ESbNT1LLkOfonsPyywcW1IwFCqfJSK5uMWqjS1ntiZy03ioitDuOX/OSdo6h
pgHSPSrd2yJi06aNn5MhTPx5y2RB4CF9Vx92yO5Eg89C2mxrWFCkVoaLDQaY02fo
IVUbd5bgb9hIvM17MCLbA23rBqH5dh+Ti3DcW8UVynNf0smarU5c8Oh80pmTcegF
6wsUYvzYQZ9OHC8p8q7pF1vFUt9RKQT0AwXkGRXpH0E2NueMpWIbaf/KxffflK3n
ByflOhNbeciosVkE1VG0ssmFvQLuDvJrtpjIu5bXu3k2w42J4EAgKCy8tmQAdhhZ
WLFXoiz1TePaxryJ7x1LIKXXLhHrztpJo6E16SGWWLGSLK/j0uLjIIbNobIiaQe/
1TxLedC9RPI/hRQ4Ti+xme/aULgBWPv4kWCyjU8kwltCBDg9cY4yXcLlbbvidqjv
UShVj0xDAF8LafUjYu0eZf/gPDJpiwXao9Y5JzXbfmQ1h61Nwbai2WLRe6cmEjBo
xc7YqCha29Kw/RlA/nWyAhqhdSf2gr3BJ0y8VCtI6TccmhvUDyXOpbEnrEKzzZuR
tfrltpDMcGdX0Gyyi79yVa6qrFV7C01WiY/qN9cBV6+VWMWb1vZJEDKjEC9KXzlc
NhUwLRWpI2e6bIW4CF72tIPzsRlm6ASB31XGpJ5HRNfTjsPwCwINgaWFrIvRcRMk
/8S0Zv7X+b9x863ECwNZSPxhiuK96BsAUV2+GcVmu/WLjNNTR9rFWU4Dqo2sLZHZ
Ra501065bWjJnXkfd3LKvqIW0NqBMTGEL1R1wQOVv/efZSl6owsXrHzDufSFdrDY
+tniKiKY9WZ9rs1jtogg1bCpkUUKI4PNd0vPtPSv9lZMGggtnJzMBHZIr6W7/oqW
F810PUWCRHaZ5vcev6SE+2deRqsDjOdq/m2DVg/o6ZcgxQ6FdnzdYHZq1AvoSYTc
1zg7Is0CO0ogbVXpdfciFVbILj+gIMTj3aZxMnhp5eK3GQJxJK2cCgZ7x1b5uyBv
NOHnQCeyti+nG8cFI0LfrQm4OsD3oqGzoiA0BqVE6SdsBrXij1Q1pD+LOqg2uqH2
9hvflt8y4BjUfCUorSreivvWYxraJCsbo8QVTEm9X6Ou4em8wIfRCqCjGsHDVWgd
t6fM/tIZj/7gr0N7izEQFCpxGBVsx9pBXuHWj3UvDTdgg2C8fThCoZB9qhgy3Z38
9QTy4mTVKGmS11pqd3ztDi7CnCOZOF/AFkIhQlRsflc51sIEDjxjDr66qfm9z6Ie
FQkS57cvSa7SgsznJgZ29FMpwKPufzfh3kBHX9jGddnT2znYEimqqBhd9FCOU+4x
J2SMPV9HiJVEWPUqOXFCNIatK90fZeqYRnOuRf+vLIFOWLjrA52Lw7CtGYwmNezc
K59sIqu7IBRaC1+yAtSzeic1et6y/Mli2Itj2eVxzWLhuzwfujj+GV8q/ktFda0W
GIInD94dQYXdhPCzsq9RtaEclx6VTxZsxi90taose19OdDYnAg2DlmsCcV91zn6y
HNpBb1zjzQTem4c4MweqKNQYRYYikmkJRCjclBfsNx4aPDAoPM5v95H6+clnra/S
Gnn7cxvVF6CRl8U0mZGKuPiiBMfUyblMmXFpJHS+1Gs6V0Rg7ExaW0Q6PXPx126R
Kj6ELkERKF0S1DwRG9dU8inca9qHckc2sT6ufxiJa11Mc4N2HxNk+eqy5cPR2K6l
0xvVqMkWUqSWMM3WR7HIMpm/5lwPrwRnMJPi9sjFqYadpuejWvB9L0iK3xwoGESC
dmPzSDx4dPHcSo5N9KH8ZGxjVQYN1qoFmE5seTWrXeIKb+2ViTMbdUvaJ6mpTXAa
8fcIzoavaPBFUR8ZYzTlyO9pvmbAg+3hgYZabFe+nBg9UJ0xqD/F4GDsyyQZ2Ppa
g9vGNSYDng+5B3VhSlYiN5izsaqndPCDq+R3oXDDJ9pYI3N/smhcu6pBlWVkoN7z
EQSmS5Ko60XXRumf5KS+qA4ht35N2W5654rXwNE9o3BBAFEP6hQfhd99jPT4mGzA
LqaTcObGCvHbRgUBA1miChi23tNY8Va+z/AIII7m5oV8RMIoTY+dP2v3OEIvSNc1
Pp6AKRR3VAkX/pYbP3aq1ZZ3264vcJFr+hKJvPa1Xof4aQ+ac1Gch794maMQTuAg
mH9/Ok4jxNwCT1fOpsMX1hU5+dxqKI00aKVrH3rblHjkSNA07l2dDvn+kGKq2BDE
9tCxQA6y55T8tIfUdVSJXW7G4KNEEI45XFvfFpERtlXpKfRBV4SZ2/6/i8Vwglya
pao50EAEi8FM2H5/LJGhpU3QKv+QpPnLZ5RLYys2XPbzIgUa9xDIzhmbtum1xnql
78LI5xIGaOhl+i1Z134d4Ob4VaF+5BlEYMC4cqIXG7gkVMetw5wqSSiCjU/cZIEH
Zia3TqVZ/xwImxHAdBx0eJbWopSJNdPNK8Hm6MUxHH0VvulQYsMh77VXGxvgA/h7
ga8SJ6mbjV+9NHQd+cOK31slIlhPNrprRCTZYouqX65V6bdRGfSYQEuflQQmceYb
RWS05dLu3e8BsKiWIQcmNsjQ/6reJQLwtgg0zcyT1WOzAD7XNsnyajfw+CgEiwHO
eW5b34c3DrHWUzpPKuGumix+sz1U7xRJi1yKV4towR0gOOvTQcJ3L4t5z/2FRmCa
Z9mZjWFLnkagdnNDx1xcAU8qFCpNVFyhps8zez3b1Lpq4zCH5oAJLjg9nMC3jpnU
NCIIVlmq4RD/1MFLqiFSroGLe/ebarlgOOLVC0TWYkuAN8vaji4iAr3h/Q9u2v9v
INGpM9UxgPnDtwSmZtXcHewk7Mz4uVaXNkeivSj8jxpXjg0IhbiqS1yI3mJDHJZt
x8z/fBhBS3tWcfyhpOlfyF1Cu8gEYbW/EHRj5801QzfAZvKjNG+yxbT8HSXY9VF/
imimDTNPP0EFmEk8aTysZPUqlqp1F9XEJ17qY+Otd4nSWT9W31qnCIepFp1+zNIO
I3TtvEyTkzwC4ACUFj6OdtK957jbpyB8BGA6AI24Zyo5xN/xIjyegryxwKyjkTTS
ivSze3ijUYQREQD6/ydgDlwCPYF2x3w7SJk3LeSpWzjCgkhHxSjT11lwM5FZhkor
QV1uqRa7vdKSmj2d7swylz63ItfuhxU9IRN46CwGAfmw643W/JCoNkliWrOWqu18
+HEIBRKhTWEAQIfm+UXk63ken66L4ZLRWhK0IyLcFUVodJizLbP/nttSMrOMeNLh
6iVHxC6r1mzUQq0r+4FOfy0O60yhoFyKD+IHtF/whEyhdvlSmMcKeemRPUYwYAJZ
5VlHImoarS4j2o7WXox3RsADYG0uLRt89XoKCFuLh/hWeUXqH/CENLrFry6nOcXY
1jIdOwN+oiTHJeOm2Qttp+pkgDzsXlH0hdxSSDHkqGYQMtiA1TLhlEvGnaVRtZjs
PT6nuyHf9RCVsuCm80TtCV8FSmrHxfPC3TzvQFFv8l7CnbRVUKL9Yh+PiZdRf3nY
c6Xww8AyynA8jLJVh775UgqVUMV+c6lctYYtvQjGv1VpSvZSSU8aE1PRBSsSoVYz
U/R8lDsEdqiPUDGZsDnvI4oCqno8VDmI4Waug9o1KOeBO/DEG4zbUbpGTKgFQ7aR
hPfblYf+AZ0/57lPEtMmoZ6dsu/45LQEpRpnjMrzdpWxJbvnCSYgxUbHt7pMyR8l
AOOEecRRf5cK43ZW5dilvbUUzJOBJ9RTDM/dr8ijL0K3vIXM+yaB+uO1FMjVB4E+
fqiqGEOADrvvIzeC3cNmrtpE7+OXFtwKoI1xZMy6AHQZjWFXLQoprgKk1RzzPkQM
f7I4eZHlOREl66nks/CERlEXo2N9AtmZhfda7AeBpq0Evfy/9lF7qutaBVNMdFAy
g32smPa/3qcqtPzIHFUe5IHZPYKEsBdF6tMrc5M9ITFQfA2C3LVlBZ8yMvlyyq3X
JDL0EpFer9us9iHWocjwO7s6oMKeSc+AZx9/9bWgVsVim99Mq4CNjVYVajSXcscF
9y0jRqJeBHifnnXDz/RnOA4njceDJj0MzD1UeDVWXruYc3NwG3Q9uxuC8p2trUyE
41SKjKTatGCTyXAvWQUlNc8R1ZPUmtGizZnXTNREIb/gi62D5wmpDquoPVfqd7kl
6IP/U+nth5G1AOqIclQzaRy3cdSIfARxcNPoKZot3c2CMSXl/UzP77LCI18FK4ra
xcrVN2NPSaIgj50LXUfp4yno9fDGSg2MEDLzObZWG+YUAyxtM2oin7dTPKhShGwc
6i+JDhyv0oYQed5dz4YmwLRv+bwyKiV6CmU553a7X8frGysUbAsYyB2UyJEBP75j
jaZLNmGzZulImSL6oZKHw3eAbYZTZnn1Y69X7qtyJaW4UGlfPEea2FiUrfYLYfz6
97ag+KcPbkylLEf1LUr7kEMei6VI1zPZp7y3yRyFjAVXMUd6m5FEfCBtpljcUOiF
vz+RdYc/KNZ+MYzYolBBSxnXyqXJrGtO835TWY/8kuw2Ris7QfqeAZnZ4CiB9kpj
u7r3LuuB/loTDAJ3RzN6if5AZY0oF8cNdI7BTKvLgIUpO5sp3vsWR4E6wIozQ5Vw
KvFn2uj90RbVGbh4gVRyuj/IBW1kPoQ4zmQVjCC/I0rurzm5sJgQInE3cE6EkkHG
Se/erf+ssOot1vXy6R8H3KaxxMH06K4KB7ODYPtkX9QJOwMdeNGlad2PhmiDpaE/
MW9v1TdCm+gVYM8rx9mzpUSd7kTzx0ioN4qiC6d/I4syu006KpJ306tod8hbE2rJ
4vXJIogP6UjrJt8CE8Py5mN3N27Yf7dtPZbUnYj3EGvL7E1lLsXx2esws2IrENhT
65lCrCYXjK2i5ShXLDvK9eSTQNcvVBzVXoG9kidZDXub9FTAiOM02qKqzNX2kJhk
+d3YK8RSzB1Ue38YGywj5mpr/zOY5hD2/+P6VVCNNDnZovgag/eSRU8WU6QCM6qf
/fKF4+OGxn1jO3PJjzhsmuiIJcjp9a744ng6VBiRc/hj0usnmlSevvSHVj9woNRI
afAbHQz0hJ8yD41rrU2Z1yaCR9htsuB/rOiM/LNWlSFCsXzte5AB1pej0bY/dZ8g
Q6a91PlFDyLknCpxEnlqCip7Qxx9TNRaFasb79jhcom6H4rg5TcART+uohhv6nGD
B799s6oVbZg8rqb+wu72M+EXNxdAAN3wTGUrHq2vTLCIeg/hHw8tA0Ld1HAEem/M
lBpyN3L8fiyc+nScGB51rv++v0aysa0C18DF5g5JMK5WMhIl4ZMp4eP/a/day/MG
whiynEh8gZagxNdfbgYb0EnemWSUpoY2Bu0B1DwdWIBZBBWn401JmDJZzZwlilME
CytEY1sl15HxSjg9PVlaPe2Y6YNP8Ulr1ot8EdY+/53JUaNRwMjm5MnEuT7PlP1a
AaDUkcNDNrtONaT4Zo3BGvjzkm7y986iabjJZhqHCzoWlbGQdN2UqHIiI/QEo/Ha
Ju15i4brtbrrjj+PS/HpHmrgdWwL1SWFl+d5CTcoced9ZrLQJrQ37Y9xmCcTQIiY
TjGBg3CMFFaj9IdWi+oboKxque82RCx4BzXq2DH6pzttI5YLpwxwdUqP+28ooEha
GHVQhOVafIuLx6KRrECytEpVSScnFfn6lv62RxToIyeuDyPRhtzUH+8739u7nfYT
7iFDmCsO6MOG7zIKdZB7QGjb1BvJZVTGYIC5SbFRIf0eU4LPmcALdyVR1S0yi/cA
0ixN5qOuMV5ZFi5d4FEu4rzXszt3fClcTNU/W0ZHChXHOXEngIRlA3CPneuKtGiS
0zDrvOWZW3I39ks3NSJ6SvUbsTrMYR0WwQEyJ6ADbJoaeA6vd/d0xDIsTqc3bSyG
JbIMSXXbI8ePWPurwkJ4Y3YCH6o1RG58pDzpmlMe/M0Oe8+v2vl6jCeFsM42+7lZ
YpmIWhMlzLtXX5++QD5E4S1b6F/sDnzHfQNopTRNpXhKsvRuz8iM1+w9bavK5j9l
2JodA3nrfSIyUUSG+KRNq/DWXlaaMg4nHsj+vstTgu530bY7XGPo6S/kNjJUcIYX
32rUfdJmFcK2lQJ871XOUg85ADd5gx1FVhVC9FG1HhToVzUYERqdes0DJuU1QtA+
6pG8gdS6r36CBsJnE1hr71vkbCkYeGKO3DaJXcmKSMDw2BlsS//KJuc3FyJtzGQI
0Oc+lRzzIV0J05YGdIPPMGqSjTK0imGquZtS93HDzbs8fXm/XoD7ac9RFywMm+XL
B2oYQ/5io34Tn+0x534LJJgzSq96wmPWocEZmL9fBAWGwy1nTrRo4e89vCr+iwaE
xjAnaRC1yYkbztMmfz7eUTKnr4qy66IhznjYEPmzROntJ78hC0DW3zKIE8SLofcW
8rxcQnGCkEEg17pZH6pOhfPpBEbH9zFH8wm3xpqNySFu1P7FAt/Ev5NCVwaWICYR
V6RSUt986n99aJBdR+6OsYAo0j/uKtNIeuFl9O8djv7BgDZUQA6WZeAOIau3FSek
iieHCB2jGXABJDdlaZcd7ev+5LCvX1F1S0GEa8ay6SUml+QZhvRMXwvIEsVHVHmu
gIgIErHprRBCQo6MHNnF8SUH0L1Ukg3rD5RnM8Xau1r05V+5x4S3XqX2Ha35yMQO
j7d0CZY5y6yr8cSQjdNNQxeP7OEGAh5zmAD+lF4eA4U0SwsE+A0HSH0wAiGg2iWD
UAFa+VBuPRS9fMeguKDmyzAMkq4cWuC3M2MCcj9Mc/77FYcQSoeq+FbQaMR+U+nK
Wxkop82UV1cQwOWPbthaxKbUezcg9ho/RbGVZfUnD1xpOFmVVWrlX7/zMbt8GqoS
78uiuMVETBdHTHOpjuo2f1tRbN0h0na7TDqOs+GCjUv5ylu8Yq399M++kqYeWC0t
7RdHp5lAbDO0KwFIpZX459weIXdBKCYze8q5NFJUCkUwyGkCS4VFIEU5hNCs9TOw
FFONY5lzG/ypUQSNzb5zUv0iFbW7yBlRxzEIUu7FxSeYa36hMEcfj+8uzE1FTa1m
Yxq9/BlicgEO/72imFX22LIHOrgnxa77zlsI3u2yKP3RT/wS5B0fvXJXXi4bs7Mn
19v/VX7KFEJxQJAiY7r706AUENQFwPtmLwGeWaKQKpuUdHoI+4Nxf1TsT55W/fWV
UuTFVL+vHYQB5HqbXJHY8rhji7W9JaBVboB6uerKYtMrSCJN2ptMw2H2hAyR93Sa
yMEX4Ay3lMcJjD3Xrw3K2rOjOWYnoaTbk7VZrZMhz/8McECEjRmbis5jVmlkYo+I
b7CSGI69jJ9mZoSJBAf+NCAR/5yjPXZzq54RfZmXCuUUSFFQ6ayZIUQrPoZVZMQ1
M0ZM8xQOG4mCY6IaOiWPPLqfDWZ78+AiVdDNcJHnRIREj2i0P55DLFX88cUuFmsX
MJ9hkvBv8K0XNByReXBcfBzurdhhGg4071uqFMT8xhy6ckEHNRYl5EGhrf2l1nFU
6B6e/kK5vWwybi7cHQhpRPrhw9+xY07Q6gYimbi94EberTMCPiE97iyt1kbVAikg
LW7J1En8QAAeQyenOVZ0SYbptKt+pEzIU4JCTP81+/FQ7fth8E+tGUNZyfvo5jU1
IotJ8EbiM7i0r84nlcIL5LfEcB7k5CFN9FCwO0bxDahVBV/vvbsp9J4/W4IUyxMv
pDPgRSP1qyc80SKjwbiU39TRM74Btxd+ug3JpBk90kyww4eb61ORedTu3p39YtGj
5YZ26vp8qamWOTHsASMNBDBofGPedbR/nQjbzNBuUPzyWbN9Y+s9pNZLXt23HJzt
AdNNKjgQtAY/c1/HhIjTHB9ccBmgrg65F/nGr9L5LdResJn0zh/WK8iJOe1QALrc
JDdFqwAdLwCqkVgilgtn0g1O9d6rHylvbvCQSnbbB/OucqDHskzxnoEXpeIog8NG
Wp537lbDZv3OVlT0/W2L4r5YkSEyWNYFhwKp9r042jYt17hmi88PFiqtLSPuUw9r
n9ydMEbTYOQ8X2To4Fo6Gai5AYNl//qIwZhQNMcrZXztaCUPyKiPUUOvaS9xj0Ke
1m7droZ1XbA9d+QZl+f1ObOHWcANHDTSJzL+sGL+UcinxD8nkcCGsqyi0nAVK+44
Kz9nGh8tMj2sldy0TbdBMreZ9s4eNTNYtsmbQhvA0n2qysyfF98QoO0HbxJeZvds
0Xx1jebCA1R1GXsrlQqpFcLrYRllAqVsOggx9+jjMkANw4C6P2i2IyN5DR8mVPNs
rR1vqXVuq4DUfAwEnaRhXSW9PJUPgLY5XGzZPULW5kHr5qn/LNdbbkEKOTrPEy/y
7qh4tMhjV8z49/aVGhJ1+9p5KJtws/pdSmS2LvErJpduKuL7SsFFfDUqgj2+vWPR
uhxvAz0srR+hktW6EBj9Zrw45syPuwlVzQfM6BQsgXgzKFRcm+iy3FmNAIOAyjSb
F8NefNRJNQ34nTilI/qGFQ6PVgc4n9rRqI1aYKx99XsBcQsVMf+H+DycuxAemQUM
r9IUujBh3dy7RpRuevOOIHOagnkwOK/fIUqjbs5JOnfxpSsWkQIvC9F1umBWJjnq
p0G8/PKs0cgBxKDJaC1xc9OW8uGUskDb4MLyhKpZZHe3jI2V8vKTVvkVchTS6wGh
y6jyNGkpipb3Z2frYyz4fF2ukFHpU/txyKHZ1EBNkdpy6AtjGAlDjH25SSw3x+x1
5NtDzu2gHgjR78EZby+FZVoIV3hz3XADIGDkYP8BteZWXn47EZimyLWIa2bJzIKP
Gl7zwBLjYYKd8VzUXZOeNzIUbCSZjYvAqyUCDim3d4/AX/AVEVCl94za9pcw17MM
SoUy+Qh76PEeW/lbI2koHLufgo59uOj4VC2+m4u5q5vTpUgv/ptid/6hdhbLPjAM
5gCkYyki0z+Cl5lVucltsdFK9OM1ErO6uedA1aDyt4ilR9fFZrDDKUjZq/ja/96n
yq83GmxorExb0MXFTD6kqwCcGHqh3aiPj7D+elSm4wVsdXXgPD6Mb2RZNmBAth3s
EFEW3Z/kuna8pRLRDOUEUsK/NHU/t6HWfqX0+BtwbkwlXWhzH7bOmGgx8O6GZden
9a1bBC/NAXucU8JDW0aHn5/g4vcoK877rMkPDos7oWgJCKqBhFnvXrsy6apayFYe
i4mKKuRdJV0CyQuC++gaEVNVoeJaETx8dvVHdqbM72FtJ6XYfLHTelT1utOdJwha
vX+g+1JvyPh0K9/nQ+AyidnhTsHerGGDSjmBUgAM9GKMVCOOlk6WcjyVX82bJgaQ
C7KgAazw+H2Qed20hZvHxTKZyesbZYvW5jP+ASRB6DRNxKgA3wje9tw+e+3Fuymi
1cPhio5x6eLO/Ycp6kw5JS1mVyMPve32Z65H5oU9lpkFK2A79TDZbfr79aR5Q4dz
ix/Ek7Q3obi4Uma2+DM5dqdFptfygU7Be6wKTndomenUrA5TxJFaJPB43wwsw8E0
iG+9bWduvGGGFg1Cg79BILDZoL6CVbtOYQRrnpAgAftawlv6hd35BlEs7yKvc1pj
RXrmYCwlVVAHhKF0OlV+Aj8f80ImBMuh1qPG3bs2FRrs4APebP0nz9jSXGeu55lt
DCwexLxhTKW0+S1nt/rRX9hP9SUZsFtS+LxH73bXC9GLCyGNIXpOG0LFd7xnaYQY
kLzLRU8pmndYkTFG4rj+rtpC8runXlXekaaGO97FaZzH4eEw+pc5GoTP88A6JcF7
36u3NKgxwzCIm9bXF9IIZQeOtzmcIYe/ZYFkVfdfNRgYnRhgfXcvUEHk5KlzKTqE
MUl2v7D3m+AjrELS9cm3iSPcloKIKHasyaxMSCpX/UM5/6woFcZD1FvaZpXzo4Pp
CBqa4O8am4HKrESXSocsD6S7RLrlqqDQu4dc52ohLdHFpRvmp0sFhh0foBiN/fI0
E+nVL7WqAhjsZQXQgh3a4Kj0SSQtxEdm5aFxOKCzrw9jXeFuHUn6xIQxAHK5pY0N
Q1McF7Bejk7j5Kg8baz0NDksyZzgVg07CfJCjTpt/qgqPcyqsY1ECBN+VlLWxGPO
59vpkIfDdqzyPBm0IZRdkLPzJ/Emx+vT/c8vXLSWY1nVkWJmq/zjJWfFIsJ0t+Cm
Cr40umcku0r5JQGjj3AGwL1UkFEJhGw1fXD8SSNRiHRSicyLzhD66n/w+u5abqJ6
10ApRLuM467a7TXH1VlpIh0m723VNnPXGZX/2M75sebLN9j8JM/49LGEbnVFeTa+
bzfyX4WIZ0EpwrN9p4NJMBxVv2VWBLostkTnd9A9p1vWwXUVSYIgUsOSxXLphBvq
FiljFY+VQldAFlOhSTETaGLokGGkgO3gZiitjXRz1w/yS+ZOq7zAXKj0lOK3nVOk
qmXxR0hOO9cy9FxOVpl2pRqRF53Vdhu4KZSgkXTWGc18gHVtzl4baWe9Ke3IF9bV
QJ1kXZPRxfcdfi30U1IimqusZTCXmM0wtpNdEYwcbNWSLxHjSZ4iZXexTsEHAaRm
xx+lxFV6xerslIKwoaqA6g15rP5+qz7r9IfVQy+S/Uj55Yyoo8J/k1SfZuvlsPwM
5yKyv3L2oLwcogtonikt5mwDJLv0ng8HLA0yFn7pz56ffUp3HJc8VpseniDaVwXS
Vjp2DGlK4QQd3Rtx35QVKeWUtB3dRpekGHFjhyfiYmsO/YcdELSJ+0xkkYvGswM2
T9/zvmxgiLWRLL7YPqxqKVatC3l9SsdqVfmYU/ZKVzwiVllYUZlUIDHHAtwmWRug
qk9VRBKUZBlVezK26lHPT7csINzdl/8ylvy7gT3rxUNro1SzYuNDEz6oY4KL5wFt
ZroSR745oS/gxK05wq8AgxZMMtSVdZi3YFYtwkt+H1PvzU0DrdIE7a8dC8/0rYZo
Hx8CCxE5eOqV68oO8cvaaOG6hb+z5cgYeSkuU/l9ZnFIpk0e9+SSKezZUktEUbPu
oe2oLA63YRh6I0DwHLHEw3Zhe64pcCIR+vHQNvgtpM3vKr1JcCGJ9ZRDevoqUWhc
4myNb3munGH3zKMYecEjoFj1XMeT7kC8nq/opl5CAcFc4tVwhwJQ4l5BFY4WVJo6
asPPyTtHVsV+SkAkoQDZ/QvWvUl50bH6sURWxvRUJZia+ISM/o1ekqukqoM698ew
FSJ4W6WYl2YxLAKi6uapugx+kwdkM3eKBGjrTUpN9vryxQe9AslvK/gYOmgYBzWv
UyYlLT581lbooLOoEZnRN7UnVafgwxqET4g/0Ye/YGsGnJyiWiIVvZ839sirBI3u
qFkBXPLpkZOicci+EixGEH9GV+JalqA0iAIiZbRMLVy4FDUGmsP3r4vYLTXYhzGd
eaY7WXi+Vy00zUfyYgub6GZvTQ93n8m4WdWw8aUG4bwF73bLBJylBX98eLcl9Dky
fgdYUikVphhBmr0nHyzZegzOt7erFb4JN2GQRR8K+bakTbZSTVaP7CNgAr5ssexg
hIr0GjbmUyWXJA4u8cDopkLwWFnZTwN55abz8Igs8cjAbHU5aPQA0dNA1rDWTixA
FBp0vJrxRGaJWe7Jcde3cL+9lrq+G0E2yVbtw8GLSkTOi5z8fKX5xMikt4cPCjE2
zNVvwus8py2w5q5G7Le9xmgv+AvNQmVz6xOaY4CSH1CbVbMvSPFnPQFwS8FK3hEY
4R5KKPbJX8jbEIAbL3C07KIZZ6LHJkcIO4zOlZKvpZxDEOahv+JbFfvTb5kHDEDu
GrQs/tO+r5kuD1fKJ3SzxbSqNZgpIqRM2CJ3Ev9tuGyjEuRAVsNDxMa16RTQf3QJ
EkMJz4eNOLQgLADBNLBFxNtrMwATwGB4hOkI5szUk0QgdSOu24zba+EEVGsErfJ2
A80HLieopGgzLTMvUU+2J8TFSruNR/kcDu92VEysMFaRurp8egfa1eswkQ1dKfYZ
bw/2nWAbKQgXtOubroE0AwvYO36yaTmOE9Zik7d2AmAgpbHUJwum7v2Knnq4wBLo
CDrl1IQOhvlbR9WYYH4qFCLfmxUo0RkhZFr0pEYiAiD5yd6Ga/4GFBchRHshbP7Z
bAk7JS2MVtMMpqOtt3ykhc9YCWA85kOfrPW3OHcP+Rsnty35rbKk2LOQEJemxDnL
j2JD1nNVb9eBGh1DtrdtmXFsDae2roQBTWJPaR66X+UPP9DYqqie+oQAy8JtbiQy
Y/H9BMhWHfI8pxC98qYGYartB2iLlIb97shl+6J97Ovp2XUwlEImKDBYiuRHjss5
RaoU22mzeUsv8yCgJhght82AhmnzH/rp5yuif6FwBT0dAIxsjRgrlZwPjhjH12J9
uta4r880G/a6KIJzl2lbc0jW/lZ0kz4JpDoSR6/AUevTKaoVDuH/1qtcNr91FB9S
XryWfecYPrFCUSBTNrDuveAlxNBL722XscEVH9q4TkAT94Nf5dj+q0m11guOOl4d
ag/apHB5OUkfwlherPmTPe0SbUKrF6BdfO5wTbYeybbbaata1tKYoIoGxrS9GqR0
q55wGIP8w5FA98B2nzIeAXeSj6nJhqhIr1OGd1CQvZVcw7v1aiIUxXdtOW6whWts
uj/tsjPerMZ47kBT6cNr4G6oVsrYedtd3xnlkEDCKKYBhokAUwN4TR5UOYjXNbwS
PI0fWyKAVLBTuMWYkNj39FtQ5wrVlN/ekd0Fcz1ojVfxWAzBWw+Y6abJHIAxFG/S
njEYkSDCn22EkQRaJGVML8+LdEOD8ccGr3WhhmEUUySuUE9kZBF7TJCHWarsqJdE
1/jM6Z0ChsaiqHMTwkTH4x/YIBuZyDnANykA+rZwZ8tpvz/AiStLqphnGHb1KFLz
nS1bQY/149bS1B9H1wfOuXSjqRM8DtbLh1rbfFDxx15ISRec9hzkUvl9B22/7jXW
ZMIcATjgvz4o2VEI2m1xC9jAmPIXi8RIVjsNZ7gUpylYM1Cbl7a3LWZSNSiTBiK5
WBbc8L7M5dzIU0oA++9Vk4Uqxqoex2JBtl0fuRiFUTfnmeoXOMDz6OMq+361/G4Q
VUd1Wb2Y30weng9Lj7VQFEc2ZjHZyTYJz/3eJ503n3Un4CfPRBoIFgdKv9vP5MFq
+KrImfFlS9ZhLVBKD3CnHyjbxiroitrVrprcwv1i5+DSGwsLRmNlfxXtKi+/eMwQ
o+XH0AmjvRKMS4CwJydFQ58ePPRuLg3O2vGOE1xhYrH6kUz7J73JkRUHlCf7NAQZ
P+cfdGPapg0AYS8PJPJn2+2cX+9dGPZxUVPGlXs3rSQDGJd96KYR64EPSMQ3YGcy
90uamd7NXR40742VPZtTTTxToPhaKVqEUe+Zi25SW1XjFzTdcvmOJx1i7vcjU2kp
ij5bYh+IUQIml76HRlRfwmvHgil7KbgbrJy2SBcdfUpQ+3rh0t2Yq26KCN2icQex
xvzTwiC+owWrglvkNDNFNCPbyse+csMusXnpcT4Dda6TOMT+mZyJ99F4MhnaQOyg
pRYNJnO4qRwa9M8PNID8PfZYM6beW6C0bN4fcRlxV7f6VkrMz7bGCt5l4xUcs3Ze
1A0htxqm0a0+Y729xBi9Zlstgc45ca9jJw2m7vkjF/9gyabI1mhM3m/3q92OEgHS
RLVIdX/Sf45XAo3Ee8ZDHmyxZL2RHM937E5USyI3GOwOGUmjC8kddwDWaO7Sb5tn
g5d5uhDV8Dv1kMQOo1k220JomPUW1U0EuDG1Jn0mQXumYRAC/eE+KeUFZN80g9VO
0QVw2JTFUazvtN5ZOPvOhERj/TzhE36IC37kSujKYJT/U4YzvXAXSQlm6MM7W8RR
feUv7dFFwp+lM666F1FdGqgB6+FCAwBQ2yGsFKmeQRFv7CeOEwwH7Q3huMj9OVcc
BPoKmEkcJzct7NqW/FIUCqjvCSKlIcPG5uW891hxXcUnvvYSmXsIhY0AQQMHTnw5
S/8XZTA8kVLK0I5CjgJ/ZNqZjvex40kf2HnZVRFTsFkxc0OcFHdNO5HiEzcJd6Xb
MBwQLfWbRynUOfRoIkWAznEv/PjSojoUhVQmO/Ipv/Jx0snZvidYpE/JJdCWNfE6
dldUBhWF8JPh4itpQrQtxr8ItuDehJEf5StMdEh4fFUwwOz6Ry2IJBysvCxl712l
HcOr3DIf+jNpeRNKeTtylvOYUWwkNWptufHvBnFDN2Q2Q3/E8ppIZyCZvMi301UU
xv80+4E4pMbNJnfirruamHJx1Zc0WPzOQbQNicqBoblJ2wQs5gVQWd1N/nLGq+Ap
Dze/e/l6aTfjfJGLfczOcN5tJAG2X2EK7ogfdksTw5c+1N8CLMn3ywZIkMgz1il1
N4nwqO0xGrBlMghetbxmlKmoz1OoG0lgivtWXCB4XZJP1XPP7z47b/+tAVjnWlcX
66AY7wJUTM6RydtsSyklybXX8HO+dI5czj8miY4s4iWO+aVrnNTRadiHnf/mctqn
TCrxfNlTrkyw/y7AR9k53+J0d1wtxBO5eBA4qhdDM7EctC0zkyGznyFbRkPoIdJC
WZQqm2GUrOXxcUVQJQkhv1+/igO44fBV8XPj73jfM9yI5ZqwsjMGoBCPFPaGgB8u
ZxRgYwRE6DdCW+PExQdvEnEOXqCPfzib4Ebry3eWRYeCMB7+pQb6o1fh7gfkEUXb
lNVnNxJXi9h/mvKByplD85jEFPsmcZVXhAo6BdEEQquwOFhG+V28eYxUjp1sxXte
Ua79arDE91xoNQtFDirRFHc3ca5Gfzk8tSwLYP5f/N7m+meWDcZuW20kiBkxhi3Y
y3CN7M/66tu6X/cDYkw+TOh+Ce5fxVxh4gOOdQ9uGGfAPalhm+YmNVzA9tE1KnF/
JWf+IXzCt0fd9uNmh7kxk1mEJcvc6WLYzGAeqUTs2HvKptOj72BUZPsLqdW3Dlma
TOskXaUHfbeHsRMkPp/xomIAe65gQgeU+7M8Xwy9wiho38fueHZm2srBDpgOjY42
hyVX3gyI3s/hsJex6z3cTTgM077Z2wlJYmz/6XdBAnMD13p7WaTykIdXHSttWmtU
9u/OnZBlgADGaYBr0KUqDfQHLBCdcLj11KjptcZfOinGqIrfPTUa5NXvsGeIrk7D
0VaETzOrPMgkZZybFuAcIW6nhjxcpIRkxvhs/PUes1KjRUKo8xof3mPTPPGX/YKJ
32U8ATpx45bsVgnwS+V1xbxJELhOBKDCHSoxzmr7cW9SY+oMH9oLRJmXdrJtwjpa
akzLKDhD6zgW+w1fAuEDjhROeAC3EO9r+dV+fTkjXNRMFu2jqXZdn4JPWGq6uLjM
AdABADVvnf7qY9N8NPz2P4i62Lie8BEi1yJdgrKs3+eTXhfBSd5cTLBFNZdV6GLm
/q6GNc4b+oeOFb9q6EaGWMIZQRoixLab+EcVuGDIvolpxTWvBnjtK5ka9velBLKM
teWAif+vr+JZEiEPR9J6qdrvLwDc3FQ0BdQM/CigqmVZz4pzigAMCWkBdcW1dwNk
SRcNEVknVkrUXvf0GYgjn/HYZotU9rLo0oOgnNOsLBx2W2YGgZwgZd6uTiD4JNhY
WXaKmKUHB1W2+dV9nhK9ZqKMF+mpVuB23riRKqysCyAVV2yvF2Ef26T8IKpuV5GI
GYEp+FUkXJ/U9sIV7LB853ErFRCaTyH/FRHzVuN29hOkeic9ZbCIp85iD1QGsDGe
bHqQ80tHkfjzji+XdOSAyavWMh36uU7rih9xVS8NisYBD/O8j6xI1p8Yt8XOsOaU
1ajsmpbFSbGMqi3Q59UjHys1rCRhoBzOkE4oo7a7AoCTcaXLTG+rTzqHZ/e108Te
itHqO2VFMbXtVplvEYRV8gVa3rgpWaeQxUBdl5GuFY8pvAyXEL7psgczrg+ySCA+
Xnq3tOn2nI42V9vr7Vtf4OTt2y+Dx6TesfWzLtHnA8ZZj7sndPQ5b4DfqCgSwpGw
Vz11lIRqRTZ+gr+6zbhdLcLk/h2SOzaR9yzrL1CUaJpciDbSexuk5qDGNSCHXS8j
vlCgQl0UL57xFAVpswz3v/4hR9/tGPsIuzidx0zw07WmeSS4ysekWZge//o1xLtl
UjCP4rL10qVPMscrmZ9eTz1zBw0Q3f5n683ampZjvDrJJ3VhoGYR0ZcsLEbzjEwq
R1DL9d2oTBVeR9fR1H+qQDDhe80+w6sW00rpMPCkfoFew+mnGcG+KiFnExkI5ZxS
p9gtammohQz3RyGWo3cqRt8BpM4hdSjb8Va6ddYJfnTlZmeR8gXHPBnfzk+Pi39d
Qyqs90EeRsXVmdIG4PPfNhJwBq5lbFoTrNyn6wc5YTRvTSdWoSDUz3HWtzpKMjc8
JjVqkBcnzuyZxoCSQ5+84SvxXKz+sSRKZT/tNTOyPuYfK3FRywzjZxjG+PvZvUEW
K/tWen+nxFdebAvWMDS+zB2oapWRP7O1e1nAijmieU31pUOW6CUCOqTA0jXZOmEN
fRqhrwe99w2cOfAhldpsvTjggxfb7kw2hMQcP8P1ezFvKF7yt4u8GZKIxsqi5x5R
cGfCieFc1zrn1fETs642THiTCqFkQuPboXAAeb+GH95psEoK751wYXe1QVl2jUAB
+W0Ot2FPXPThW9WPWmff5O4PpHOlIONJ4c1TWXYkOL16+Bx8DfOQL4qIG/y6d+Dr
pB8LQDdYeVJ9otfXsNK7sXhTtIMIGsOEIFY9RUhG+72IfVTs2rj/105+wtmdaloU
EP/33KvujtsbMIwFRDUOg3I+/UnPVFTX/pbLyWHdVxaBxpFPHwUgWH5HOMlxfsuH
gFvJmGTQ6qSzTLxHlFDrTgOC7gZjZM78n4+ekoEpes5HLRCWX8ErYFCaPF1VpdY1
MRqW4oa00GPe0nS+F5DbubXO+aJrA9nSjZWhyWmfYfa4U1QwWnV0kEigr+UEM422
sylHQnW79lZDpqAjjKYv6pMHeWq/fbc6iXnjkrSAeORMGG31oKyHEK+8/hhfCMlb
ubdvo3rafyUqAAXP23bStrBd9qpaONPYRrR18yS4b638oo9PmXZZUqMViMxfRK/c
2JzQw2oSOEa4TNLDQlBwTJ02dpUiPt71k+D2mAXrRUaCeE8gIa4Pa300se8oeyAc
M0g1QOxJ4Ij5N5kj9rbbXG5axO4s0SemMV82hHZ2dakLt2reQKEeOW4bfygp5ntZ
6swTg6Tpwnb7Y+m9zaIxkrbWlMi0B0c0ojvZgS8on0wroJ0/t6U7eNTPW2prDJSI
wk5gC6EomPKL0JndM5cT+YVeyzXXO8yGFGYr+MyrVNQhYtLyh4OcZ2jnu/pX7dae
m8h1cTRapbnfB1F6jkTtK8fb9l6BeGhRhxSukOU4bUwn+8Wdxy9M5naKlasUmwzG
F6/Qm2mDuXGgmm/fZV1eZ4tQC8GwFMfgnpi/4oq+2d943N8GYu6945XNZ6Av93RF
L5jc9DHEcGyLCyTL8ETHa4IiDHWREU+uERaiCMA+8hSXD2UGFzfKs6QWdaz2qMPA
p4dQr4NeMkC9TaITwVWQoUYmiURmwFDtvtUb4I3osG5YWG+dK7uIf239xcmfAbpp
RmqRG0BZA7/eVYbYTT4rjfgiSsAvRDhz8F/Dz3hsLmqFS3SE3MlncYPCRzxHGnlh
Nv8/lXx+viyRldw5yxqWGlbXfnkQHP/UQU1lQUtPdXjgbMdu8BjQXXc8ZH85vK16
YeXhmsyn9o9sls8/V8Y5FkfuCBoDLA8LHLZkpd9UPnpIwgMJjz79ItgO/aLZoSKj
IvzlL9ci8XGeIHF37AAz1HJejaRfADe1CYu/K9E6xd4GRdVRHED/naAAEQp5rbTj
GTunNk2KfvWgVALP1ojQwUMcmei4EZwljw++0jFQ28MYkoHTNFdp81lJSfE7eCbq
hbIjEMvntKQbHAupc/LUIgVgVIQG2cjeTye7J61kL2R7ncetQ/0BIPeqx7nUJMsE
u4gM4IpJ0++nFSkp9yDdCgD644uGd+/jURRBg75hUyxanbb+SfXaEVwhpnJOtiJ9
f4F9/3l7mWAw9CLAtxayMvuhJ0KZW96pR3D2ciBla41pJX8FPpDC4mmT+Cs95vrs
EmfterBnGE5WW5yn/OZio3ro6bn1Ulu5kM8qvQjifJWA6xJ4wPh82dJi44JQAp5l
l7FVmxRgjhu3ZaogFBKr4o5ewcNPbv0Gj5eUlxp5lPF+TjahxytN6vWSEdPYrYNK
HWZLz03hdobRx1JxtZPoL2VPpz0bTq+rqOpe7n5gAN/U4aLQWCfy6LDH3daJgjam
vuURjyaVKv6L6zcmM1HHgH7jUfGjhk40ucTl/oKoqHKlGf/gdKeGV/wgpFgs9TQD
NKkdKwzvOhFOmdtRLAD8O5YctOV5eXy4hPAfJ+xevq5kuDQ2Ai4BSr80BDOB8ose
ykfKHgv0Mv//VeQwwLudnzWdl86GOl9/MdbvpqtJoyw02eSoOrMuA6PHsZrPVOyq
WUxzPMeKfKf682SlUh8v9aFKdGmLeRAQl4J25ArJSFVg/h9o5nLiAeFUWlL2CgZV
YMgNXLeItRX/WX7XttLPbzmNlgu8ngrSTDY2awdCcUwxFcc7sp/4CcUR0ZPMpYh/
VRBbS807BmTonmpOsUelWQ30FKf66Q333xzA6+LnUvctFXd5zsr4Veq55xUSiUwm
l+bd7gVxwDEaC2e/X7RZPFOIvUq4NVLo5iQDc8+Eenf67JufjKFffc8wvIZ78Sil
r0tIhBrn9HzVvQeqz3Rwo4b0Ii3iaVEyeZ1qsIXn/TGoy/dOThVfoaJ4JoJOB66B
/qOeCgWHgWCVF1GDS+NdKtg5ktxEcudDsGAPzjF5Kpx46ykcMT6OyXlfjhUYAPkz
e6PwfwPbLadmDFJchhCZamuNjCwihCUV6H3dCQN+ZX0CyaAmg6Yaa4Qji7JYISZj
avd1F/G5CIvO75o4vGp1uZLaSMS7K5lciMrtB380JS4ceUDXTrG6Gxc5cN+bWVJY
KcTGR1UG76kawf3EQ9Vvl1UPnIltB7KpNn2SCoiariA2CRYbtyROvgtZuzzeGUp+
3NDiDC6drlSuRHPvaOhd8k1C1Jilt++Hn8PNLVUjnmsDxMKTZTTse3vFGVazpFC2
3m3onJxooHqqg9IQ39ZM2K9o1H3taokow1EGdhyloNZTG92ulxq89j6R8Ho+G6lg
5UlwF8XeEBzpMe9GyQZK9V3TEFSREM4vuZ7zBkjQs5VsAbKVnVuuUJIZfYi2r3Rb
V4KfLNtbTbbMV7J0cWt3YBNKuH4lc9pgn1kAFKpVcENNMCiAbO2uua+2ZbDfjbD3
Z7Hf61j6GjXLyzBDCvNAxNs7f9Z9PrOXyLnid+20XgQ=
`pragma protect end_protected
