// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
OlzFi+Z6GWfaccS6TgMgvaU8QwovTxH2xSWMGNDW9wsA16RI6+0TmPUMoMHTn0aP4MZ8eOqwjh92
BA/1MYKPDX5aFZSzGhS4Gn3xA7Zp7hCiN3tGJCd3flah8LFJYDJcIlWhYHlnGfcSsrQVZx2Ycbgm
w94iceDMpYVNbGIib39c7icrw2aXfZM7fvRtF/f0qPIvRw6VLe5tYTe8/Lmzy4qoKP0+JjACeseB
MbCraInuPupjSP8lGtkFgwmeBodu8e3ATr+2aqVbdaAmO40QUNR0KSdNJJvQy/aSL+fxma7OrZXE
njW+eNadbWL52giNkKkRC+QiR7mVGqwDlSrZcQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
6UD2sD+Q9kiOFpi/UaQWRMpxgaNu8Vo1BrfKJofw17vtE0o+7ipVZ1WaEgFHsOgonTP1I8PKN4nh
j+Q8cazzrY6JqjzKBbq7NE1K0SE8f3FOLcTUqGwIuZY9EkxFJIed9xedMj4I2ww5r8/f9ELVsfDh
Se//E+CDhUWcQt1zZXZVqgpV1xTbTyNXuVHQJd/HJw8CP68Pz3WpA0i9rjCmwvw5uigXzktXVU1w
0ywMr5VH83kMztArIBnmIf9sqzVZCeBRj+W/KW+Z1OtRsetChxxuinGfUoDkh54B7c5Qn5RNAyCi
edmL4E86FAx45nF46GejGpC5sUJNhuc8syTsRqSuxIZCrnGd7g4p8HOSL63NiMsxoiAj58LAW+/A
gN87TK++urEO3eqUY5+EXlJX4NYYQkj6v0DKsFyAA4nGs5S3rsS2FZF/0rn0Xuz386U9Y3IQkc+i
944f9XzSRI85tcaLutDhvg0O8DoAZ/UUeM4qhMG+Jugsaj/PYtyymx/yk4T1swGmYS2Apz4anefv
gz0PRIiS8VEmHrXyiCZQ9J9W4W/6oJT1OU8kV9oC/w/TMPGp02a1mCoJMwi3gqIqXqpvJMPKVVx0
0I98uXIJSU0YHae0dsDenG9/+rIR+vx7RT206PeNFRkTGYXdFeuf++PWI+36ofZNABfUNwH9qRGQ
e7HrureNvCufj5ofKPDKslFJFf3s1xvT2pcuHOqZQnz/HqmF8wYg5sYDa1K7C/b4ewux28gmFf2D
EH9Sd2wwrayLY+Pm/8naR4LAdckAlKa4s5DxNtBm/aTrta1XrdUFDQ5TjVXNzpNFvG5xuntgotEp
FYXLL3uhQeL5j71Nzw1kZ8R20VoOhMX1Bh3YwyZ4d/c8orrclStAJkiLIWirz7FY0PiPOhqJDt+X
2KSj0LXF3kZxU6U1wBK622fbO8f/9k8S9p83qnfuFjAnXKNCEriquGuz8MKAo/oWN7LwYCvf6t1C
5/geDusRVyytLBz4YMt6M6aAcDiEtTAxK3c18O7Ns9oRMP21TlH16910KpE+3iOeJIKwu91xs1n5
4dpz/0jzpQd/PijrKnKo8QZa1Ifzr7mCA+qxmEnJLjG5DqAFVVePlazyI8m5pMEoqBwtKGOxmqGL
/3Q7X2TKUhTl/ZAcwnqfk0WLxOtSmSzHh5kvqrbJISevvrg+akOrRLR03kKYSm7v8xKsZgtDepNb
9Q1Q4EmmIfhvnTh6ANmIovBkBLH7rZAXYS8KrH/KYEP9f1IqD6t3/NA272r7tDoC3+HMX9HYi+/v
Qq1xp5kX2VuweTkiuyEcmyN8fRbMEv42T2O3GmpaqpVfxQi6tiShhRQx+66H30dL70UnPEcz7oeV
snHJcsr7uLMEbv/yX2ew5tU5QrI0Aj8fIS5a0NuuOHtm33uotZEIX5CS/WrHUPfM8CxyVpINbbCV
IPKSUI5wZROYawGTGDJPfhpnO3QgfzFE2Emtct4vsOr3gQqCnCKlNozmqDCKDZRCjCxLtUhUVll9
0muI16i0SMUG8LJGxdAunDeVlvmr5IjpY5DxN4XpE+Y3yN1xFI5Nl7sPd4+lp1KviFs1ItVi41He
ml2Rv+fZOZXJ83N2hF+08SB/7YcRkXNpEm5LdB7AUmvubxv3hiBbcWtUv82UxZjlJWRTksgQIc5h
aqGXb9VEQz1QJ6wLzGnsb9Q75owfCwdP6soOne0I7CXeTqaQNAEgdkD3lKpmFgq8wiPhjwgmgekx
jwL1qErYawO/lB9aYu0LgycSMlidNJLCpJ9+bz4hzdfxJtQqYsz+gSkPQrPi7I3MgwIM2IyT1gMn
F7VTewL+/5nuSoVyiXRimy6QP8WKxc01ZeuvY6nzuKtch6gOqakDIYb/bizpJ3oK3Tn/mXYS4VuZ
GIvHZoAox3JtQAjrDluGoh3vHIGJ0FsQhYW6CZ+SCQWnhzU+Hzfg0z0mRnIlqWlbkE0gPPFEfoab
ltAm3UUHYPyqJXbqswGL5Vz/NpJwczIlwx+V6df7xIoDwhD+tmgej7H+wqRsIbIVKPPTIrhrxiMg
FjCXEfJv6l17rE/vUw4kLiDc3q03QXaTiGhFxHQyFQA0vIj7xXcOVJLrOn4p22hLH4gGxGW9q8v+
GjBlYcGcIGvlufnVAVUROmW58uVRn1LuBzHq9vzMZgME3kW8U8UteAotvt3bIjNB/pRJwC/HmhGP
2UEXQBJWa0moYm0DXngBtIun2HmULsF/WnzsW46Yf3/cQrE/WRAzYG3mplb8jrAOrrEVZipj22y4
BIGq4KxYK4FgW8Yjh1ikrO1HpxV8wbiDVkfo1177qbcZd+SPjUoXgBwJ0HwlmT+p8nboMgdIOcG4
bzAsy99VgI7sk/S3i/35IbWJjyJIq6gKmIkAOYcDJI9OCGAGWBDnAaBUHn/ED7MnNd45jDp8DRZ5
YdusezreqnmHJu5oaN0u+eVtBqcA140Du//rZkYrAS2X9ncpCKdaxAWnvcalu1AtFi5+LF7tTtzB
1nv2HvWGtNTlUjygNcqiNyHZhm7tZkEVMimsFsWNigCC9IkCNz0tOE2CUJeyhrLhG3Rd/eymCrrr
pLhq7XKhUdVF/FY3+AzbnKCqea85kSgAljTLXsLEdkffFulWvQQ93htEmqv3TWcJmUGNYf/BZ7CA
fRMokSnTtG/g1bOdLCqmhXibScl8mHpJi8FnQ9Ubwqe0JtSdhmgyNZ5tp+vwdRKY7QK/qo/BKNPW
glLS8ONOiTSRmB/gd9IrJNRuZMfyN/+GuuWt5R7WN0teKo64E/Kecp8fI6g4nVoUe9ulZbz7D6tV
5fMWVdXCH6H+CZAM/voWCrfYxvo/zO7znYVn8LAa49c1mHWdek11nzGAtaOSEbhm2X0J9EE06uBO
50kzVDSgE84WW0OeTFxWoOJ/L1IGvQIoT4JPvfHYJ4oqKFy+LiMPhvH0opFdD5sLOdhqzlF0kW2x
b4mKx2FiYvcsiUFWriKtFwDAbbPxeVQ3cODsqMzmheUKMujv7rbOI0oZFGfsylOAd5qKwCR/F1yV
olUSsORek/ekEk9BF5QzFK3s/jBXBsQXh7ouG3fQX7EzenqmK93Nb2kapuqHzwtqRW8yaY0hMGUR
HVrTO2V6JIJyFIQxjkBeYUla9baS06WGfxzt8ZclL4gJ2CUBng03CcQgyni67GamjDyIKXZpQR5l
y8N8183KvAZXJdjyYObyqIyCs/oKTdFSQr67J9yPV8oCdvSmolHI6bAtlQ9DQ+tLuoUZrHJi5UEz
Kmnu1aya3DNq5kuHPiHQj6hiRoIhOi1RFFhBPiSXoEHumvFFUvNG40ZNDpN6fVLQr+MbUeGS43ZO
VdND1dzUslJB//jNmBZn0BhudnDJNvUkm9I+PLC/M+zjaxjxy5bGyD2H7u2iAWlvpumygdR+I5m0
czOlSga6BVBnHx0hihztOnNi0iGSLtCqEnyrNcvQyKuQllUojZDTwZKBtFb+6IRnQAv2UPQuKdYb
Ea0cyNOJpc3jrSVf3HPlHIb8Yj8lWSF0ZwFT7+QUXFY6QUs4Yf/38LL0AhKRyh34vb2kCKCuwzwf
ex5zvU+bkZ0bCDrk5y+zIZjaal+93/RJ85hXJr+qfEyQvX+vcCs36lgbTeG7PdPCh9VNlPzR/G1p
PzPr+pB7zSoZrZzCjE6noduR14cx+X4PoNbSzUC1k0Gahd3DkWFBCkVyjZlpbAd22hJq5rydPWM0
IXQX5H0VLZ7cJjBTs+gfe/Sjt+vBVDSq+IIB0SovBN45J/F5XxHmEgOLpsKc0MM9IXw9DaR7nl5e
g3uin9wxSyfjwx+xQvXZjoIUDQb7l1GktsXOf/FSprgIOfuqDegP3wvF6toa7rEXEOviZsXLqT2I
I/cQ1H13XsHHq+dXb7i6TvzBGRvR6RPOfF03LdExLGrAaIPkS+GuSRtVOk3O1uQOQSPRsYo8uYt2
byISMseaPtyNkIjYWXrDyVFQkGzvgH8N7f9kUnChiFBaJOCBNduSQadA0om6g/Jc30t05lbg8kY9
zxm7Cv9avmjOShA+4ZjHw2XzL1cJHns1DsTMYZBPDV9UlnQm6t99c8EJTLeJWs0x75oT9jc27KYD
u3b0EyH8AICEgdsgEpBHRim0Y2ohH0hXIIpXnRZS46Yv7CZ3hLctutqxtnqbRQbHd6wdgGzMB0mY
Y0mi4TBaA0V3NYeKGE4phiH+UcFBz1U7F0RmF+cIcn2C4ez4FWySeELkrnFq8M40Insz4t87DYbW
hu3Rw3OXa1jsjFAi9lpdIpenp0/aVc2g7Jsabunhs22u92BR4475z7777dBWW4T0RMJrNTWqEr8+
YjY2U6gTlmMzm0BwiFICLm4qliKL6W6d1ZFuXK5zLeT0PqiLLP0AvoGgKfxwuRtmWFED4gjz+duX
Yu8886G+qsCFesw8FJ7RHZ5h78PkSH6BsTOY5LutVvkfj5DVHEQZ+UpKyL5x9KrCmno3cF2dssdJ
XtG8Trkt+7x4QrT+IacTI0uU4k5eiCCYkXYRXAXhfrRVZofwQbDj7v7QXqFCfIfO3PNDwlJv4xXI
iITfaL1hJmIJT7kQpgGTGv3p3beuA1D3IYfpyRwl8nWkd1H4HJWliwc25ILAFF6pDqWSNG9nBYIM
yoCkOOhTTC2FJCyyz9U/ezg/XChYHJBPf/D6Y6qIl8f7vCKQ1bs7EoIsIBK2rzzZdFKlqxh47F0/
4rOoPpuTBHj2xgQBEG6GkkK09cw7LkXAbMj4u9LvVJc7iNNUIXmXZUktr108uG4yVWLfdr8/OuNg
+WEAygTbcQrdOYMWT2cSpOrBT9RH6PT3sXqyVXkgmidK22oMsksBzRpPEPymcZywSMp9FMoGuhmM
y07myfoYFtynNBIuJuiIaLQsIU8HwHgjJH9/wt8k2/EhCZ+7XOHXpyvjXO91e2qEucmlhV7KIDw1
XfByVoiw6uoUaYGJZXnorvC/Mhp2g7WleXQ5aY7NIqz/xoLr5p3RutKbpP4PkiG0wmkuS4jPMGud
P0+b7ffvElZJ6h9MmYM/jJXXmaTaUdh3qHQVUH59JmtsmNe8qQ9CETRKYpljkAv8aqYk6SkvugX9
oaqXY6zHe8FBNTPiS5OrZViY1pF+pG4pDnrcgghBHF876CUzo2b5XvaFZ26JExgxa8j0UOgI77oF
nHQoUnDOnCA+J14xSm5Nll8+c2r9ex0jGhGrNjRib29XulhGfq0KzQmSdDcbxoWbSgjns+HN4uMQ
jGtPk1Sy9yht8VvvpqOnKm45SE4bnnS+qxe2kg3NsDC5PRlis0emnZN1eTHFyvH0J8Q1JEHGsOCq
ygqRi9n/o0gredGXIOPj7dOTif7NaGgR7sCzu2O09eBncBfaFPEEdn5OUnvMf+8t1vHbDdD/0qIh
rbuF6NFXowhfeJbucfH+OvTSNcoxJzZQ/I9LfYbhnQsm7CVTlkJ68HaXHbymV5OB6XHrkEo+A4LU
1aXWb8NQNKh8KS6Ckl8usGYUpjIgH8iOJk4WpVQcxqntvPMvswyvUiTB/zVOBEIxModgo+xI6P37
nHoT2VEUEeay52HW2sAandyPjBTlV3sFzho/MH/VeXYdfaw8UeMgbJW2ACED6vcNg5+I9nh+7/1y
f5p6228K+U6GHTqfWWyAnsaMQRiqhCYrRRnotLtUvpZACQcAnMAg6wXx+F6edAlQpitdKAkgAaO0
So5BwkmddwzO2V5CTc666/f47TNMcp/IOqH1Het16KU7Mt8nd0q+H5IzCiHsL53A7MUXJCRyRX6H
e8JfuPeR5Eb6lk8UjFylSJJUI+dR9RO4Gdu1Xpr3sBrgSSU0LYI9jfSfwmsxWegaMwS6KZXqaZRz
4PmLqg0R5ZT4UwxV4Sq3tgrICMva+aNuI+fKiAtcbk5qc3M0CuqnxGU2R86E2SVecqHeXKjBk5fP
K9R9v66QwBY9yqp7+Y7r2k/+7tyLS3EASjadMWs9szODVZoqHHSUHV8B3XQlTZXZ+r880n/wPkWL
GnuYphnIIA+yanfIf7JFDt31mWpw3dP328qFxmw5V8tCNA7BHl4RP89EDGfMcF573FnHgNy7/Xqj
1MDFQhPUrhvQkeejfy8ud8vFuofW8Dew6qHOwalizo9vfIqnQ7/o7edqNgkpDRqRfq2YgUWjmgWC
zHEHEI03QNOtz8XWdIh2WZ1UDBp+kbLqXuu+P4ZrxPgz+kpQOagCssS8vf+vo1qDmfjBQppKkHtY
4MNE3lE4T3PQZxk2twX481ohFXb2VBdsYqqUM2vHbI4cHOIBcPaJZrrfkeuNnUCMeQDiq6/mcK4f
PGEWw2vNU+Bwm00zNdOsrseugLaaWwnYWbvzPdXHivbYLLT9V4W3lJb9xks89RKpLG1UjEqg1Je5
k4GDedDbmBzZ7e4I51oTNh4Xvpwx13eYCaat80kk+t6IhfPYBJE0XROYz6HLcp22FKZ1S4B7Er7l
VWi2aEaJb5mQZFWUlIXvuSDRZU8sLk4jHA7klVYNYU200QxEIwEu18rBw/gT8VW6PPQg1RtXCFs1
CUWpl29freMWsnQDj6kqbpzo6ZFUe6O639GU6dy2NueTRbuuk/bjKel0ESUGgPUF+wISEw3JleL9
xffgJugfquFGPRg3fWuwHwGBnp65tawz7yP0cV12XfYl5YqKqxuj1wC3kHmGSj3+vX5ceBc8v0op
M/pOewzICzsn/XEKDGy3gfc+sDfKr6GnqS0FeyT9+7eoNIXN7NxcUrPgO8VYvqp5yCfXtnc4VL/Q
0SbTjfjU6nfS/OGpp95WUHgj4kzMxnrVV6UPuLsnSU2ja4H9UStMTBe8C28+RhO7xEemRALichzj
CRimOd+Lz0nYb9W1lShCY2jE8Dkit1uAttSMo2XAJWv5MOFL0ffNhhQP66e2Hpr8T/7BFwRFYgiW
MvDRwoI+9K+vbYCSnIJ43gR/cqYhDe6fxZHy6VNGmLtsfOgg/h7ZHdkcDoE2uY26Cswd6bBwymMs
aHM+9R2Q48uQNxOMRSryV6zoKh2FUpcAPrhlhBfg+39sgG0lvYLIARxJ1SXF9Ou/2k7pU/aLL7Zr
x4hzEdmw1tQQk5WQn30v/a45X1Yc8U1aluBtRke3za09OoO/h4hYrRbM8n0IvQkylYaqOzFcVcO7
LNiDVLiwqPDvJX1Jvwp/EVdVoEnd+9sMJHEHiCTqZa91rzOxKK7baSf0yKkuTtAPxCCgygQ20AZW
AwJHrd7dh8aQMe22f2oRKUv5HHgD90srtuqE+vbYTqx/O66lZIOXGtVPqYdfSmJW0/aqne6NEcK+
mSSmAgcP0UFTorx5QTT3IBxa2doha/lQOgiHFnku1jQxSJbVXWbccy5IQ19CRQp9AeqJxTQ16c88
7Wj9GJFvAitpEJrAy78FBiJwi78ADuhPvT5AJvnxvLr49OtqoyiEjML1/FuUxT6L2eRz7DlrTofB
4j+a8W9M2eRT4+RSPwqhQHlYns4P0NlRa5NkpnSFmjEnyDCWDF53xUamzDNAZ6da5cPSjb663wS6
HQ9At0EwZWhEE3L2FEVxbUmh48xC+J5dMskFCQSqA1h+ZDDF3hZtp9/cZsEEZZZq4jJLbD2YoNEl
Nrgc96l97Z+PQM0dNmQlvDPW5Tou54KXuy4CRwCdUPDF5ktQUcTT+N0+ND0Lu0VzCYvHyzHuRJs3
3G7ai+Ng+olExzfgnX43NOjIh88PXbhfQhLv/vVVo/2I/kb9M+08CfZAwcmrOxtdqEzi/LwSxZ7O
IXqh3psoVxfZ9OHSZXmMtTHXvcIsPiufPOmpAiD73oBX5wb1QyueVCyESy0PAGDpa7Plk2rcIJk6
QHIRvyaDQCxICql181bTpiURsGx4wJ7jhOV94MzobiyDBtejLArS0Y8kEaEBAF+EFovOQtBqEElq
d/MDo3JBmOFkfuE4sz+d8uZWu7nrJqVUlOEF1u7FBDpO5/7OyaXMlsCb3X17URpK5YildkK2zUrZ
9rDJZY/5g5Xg5bKr3KqugrWhcOQUKxNJgrgEDKObENdoMwx0vAsa0U2HSnIggUNvOQIB3pLJ7Qlf
EAwtiTLf3Jw3JXyNltU+B1c3cNWXEVS1TYhgGGjcc/KrYb8n/RJ4Mb8NyNtGVg5WgvC4TEXZltvQ
c8TlRO/lrkZZ4WCXxZG+HJ3vTAgBJBaIhYLCYQrxByr/xAdHy9LtZ/GgJScLvc7Z6Xy7oSps1Zl3
VVyC3tSm8c158HJmzWNBerqcOvRqonOStNwVIth2hspQxTiDeegH9QzdUnk8sj1op6cklwTTEMlN
Phxq2+80nq1gfvE3+ubeBXwNajL4XaXKm9bc8f+/66hEB9YjwX/UVRzB7DUbHXPJhlmmlDBFFout
yv6JDXx5Ug0CVmrW+QppSv+rzahxQWUyTuzItmUMqIxl3SiORkRyNOhqReKZ1aOeYgcCsf+1eKBp
RK/VktirsVu54HcUkG/x4rsuAnwtirHlV9zAFYCh7dipV25IhLGQ9a7fca2X4teXpSHMpQpZ1di1
51NwovqzChgVcv7kHJes7VKCOHZb7KaoD1bawDVn3i8jdij48ycKU5k6NwYhCdAyfQbsR+JthZve
kZ3qiSSh+sG1aqbwO3/9+ofNAc6774oDk/+zTzBkSYn9bSfeVOL8SrO63dfTjI/hONkroUgAs/Hb
3FkXIvPnXWNv+CZIN/IAWEIvDNmn51IHaH1x5YsJU1v5mLcXPoic4utPhXuYmVzS16RNl5RBl2Wp
zob8+dlBlD+o2+uuiWPhJG1rM7/wyd6LUO5tXqAwSHmLrYDs+g+x8QCp/Zd6haR/rDasVFEoQ5q6
fJAeE+0DL9r+X8/olmPFHXW6PUuiqTynJw5EmKmcVKZ84DpSuxjur/0C1t124fkAnTUCbGY50Ozw
OJ+1v0+ry05GhQ+s0lnawd4gX18++m+edHNcAtpvEQX/s1poqtaxvZNLvY1EoUMCdd9FSBAgY3Ki
VSydhfMlN8C1rl0TUuLHn0UQlY9jmEWC+JkP7tT0ONOALjHCi11soOlNv0xwXIktuH1VOY4K5Jb9
h1be+G2d3nv1If6Bsh2w3Vj0f5JFEI7TY2xqe67lZIfhS4nWvcCt8Rzov663g37YtNeVYdzKIQ0p
+VEolLw8SZ3tX/EdVvdW+OpCjm5K9/kgnKdHEOPuEA2wlgoFlh788gzY7HGrqJJOi1DFqEKM4+Cn
ChRFGw+oVGAFGN5VVZerWrUiZkbR75I+3sUBrQOpCGP1rHcWrIKeOwvLsMVw4M6j4+6Z52d0qvGo
BCdD660V8WNZlXhtdJ+vuS4tdBqPVXEgck3Kuc4y+EfgttSq813OUqw1UMo+y7GdwGLr+Yi0IM0c
9ZPolBLM8loQslzzU7h9MosnJlTkWhKHbL2KdyF7IvubrAl13op/eTpNn/I5qXIdv3EpPQcvLea7
VnlM35GrgeK+YIwAehhD/xsfc6xon4vDph3fgsxLUH6tucn+BvFh3jnWIbsEGKvEp2K57ldjNlOa
XumeAne/fSvcYpfSW5KroB5fmJCuCnSWQD5b6gQhRGRxP6qnzyEGmtyAeW3K+Jc9JxBYoLBldIdX
0N8Smureh78onospZdfQlNw+dJI8VJchVv/i6Wx6iPmJdvIC8fzC8VbTnJKwjm4GhT0oZOvwefY/
73aOTQCAEQi7spfBWCM1mK1fuCTC4zv5i+TyU9+X3qBabM64sILoyr1G3sXanQqP2369k0CHq6A0
hqKZq5mpXGJBXNXGL1oR7DFARBS2o5cQ1rPcDfjbZNzZK/vI3nub52tMAE0mhPOmrVpRPV2cR5q/
zh/3S+zYihAssf5fN4KbpTnSfogGaLaJZVWiHcV2bzsGS5B2p6z3on6zyxmO1Dli8tk2UhNSRMMO
AkUcxB7YSy3mmlAn1YGp7cKiSBq5I7rhBNgyIb88qhVMpaKUUBIvk6z2tXZPk2BJdN8tXGUrPqdN
VAwJDtwFTzH9l6bI/7SiUVSouYQ3ie4jfK8seLlBjsTOPJOYzMqjZ4BxbRoQ85ldwHYqxIp0eU4e
RIaSYDYzxQm7Jhlr/V2j8M5T6ansn3K0MP7v4XB3TQ3ogf7BDvgSKj7S6drGm9U/eWyKXTUY2Jv4
IFYUUH5Kai+rNR1TYKh+9T8wwH36RuvSrMbw5szGeY2pUMKE/W1PcLz9Ev76GrsZ1NaoVNfgzCsy
jyJVhkbSXkl93pRH1FZ/6wEv9Ms8hdupTY3XAT8cx8zwtG6KxDIQRFx30fPpczXykUMwsu3jQcyJ
3URYA9XSfwbU0SRsaYkdrI2BjfM9IApFHVOIlScodPl78SVBluQ3rhQkv7uHJ7JHLLlBtVFMnbSR
D5C3ZYk9Kwec59yZ2+xIh542y84hzis0xNuYfEwaCvDosIHJlUg6upNsZyjQY/MKPQ4b/bYJsVwA
KlG+juJ/YtrwFUhzA9154jbgNg78z0yO8mRDhx076yXm+y28S7oSajedCEPr7WsXwzjETfvcv5gn
JoAS4Z0/08SsDkpRdWJHtFhgjUF74+Bp88ySEgFN76ng5LGGh5MMJLfSWMYElUcJfXfjOgsgroy8
FlxQCO/qKkSzreAZVv/5FyF8HDY1B+2cjC8dP6yYENbvYXrPv8O4xVKLZO8ijYf5YrBw9hbD7aPJ
ge8POyY3burV7XUN2qVjtJ31LMkdcyrxSu3jBY41GqCXKC8GVt3ggaZoEZxI0GKnmly2ShHHfwQx
+IKyvwZkecBlQUgO1qbBMOwK+3DSaiZix0jj0juS75w8uBUeRX/qwlvF5NJJynAj2RT4KA1kutnf
qDGOBZ5rK9oRX3j5fOcmc9z3sTtkprto+lwAjoR3jl7AykLxWjQkJfoUoK6yzPjelI0ozAKGFBOL
lpa9rccogev+JU8br35eQXnneiZ72vTygrWdU0TpOS4PaQJvHNSkBWc0eZln6VJpSqvexd+Ir6mq
JRdCccRwxLGSJDhqVuBW47lOJ5KpGqFX3JI+Rfr/X5FSkl5Xfe3hHTYKUPcHyGUJmBkKteTcUxD7
QUzhkq62gzR5olDIGmigmXdJurE/0kRk8R+rDbHrbByvMBLVHGwKZlfm0wLa4StxGH9D2Dq44orE
Ni9hzDbTanwI4RhYAhqpsNM1xMecA7odSXt42nJ0VrgicBriwFxkEIhWuFEmHtToaApUyuaU5dj1
E+dLGh4HnB7mxqqlfJYigMaGBfqVghiRWH1UfIEAwbiS2XTJyU4fkxKPPssGJMV58m8h31/RiZOP
5ZwvSKThU2kabGVx/17CHZtBPnnJ1gwkn/kvtNFw0oNsS//BIDQ/yUwWBPgYevXg70lN2bOlS6En
sb2Md1Jp843GTt+6AljAQD3VlU4q0/ixVOcdZH89pgeiFGItEv5ujfdf3snkycS91xmTZlZeVIUs
m4W041JZvLk5YORotqQczOA7MwtnBv/Zz9M/Ld0hWcD/BKxeCs+M2PCPrnfGlVGd7+LAjts1kl8v
mNgZthFL8I1eJE36mWC/Ein5QGgg3U3ysFitIfh24LE2o+jpVjD3NId5h5OLo//awK19RbPmu0aS
b4bZZ9gRTMafLcO8OqAPk3YJn0luN00G/uEE5HLZuLrf2M9Ii5vL2/KbB9JjTNaQgzLLluxsriR0
7YiF0AzM/8GZ38fe9dtZHZ0Ab/xYGJCilw1e5QV41LnZWTfr4cQoPtyL6ZQj6qXCucL66yxqXnxW
tzZztY8r1UNwyoWcpTdf3YDEbNlyjAg97dYgOFWdu8hzi6AmghHafKcZGJX9wIvoyamy2ZppwmU4
sdegOdHCE7Q7YNwna9mVqSHSPNZFnTXHdEAEOK9Yf/JpN6EAdnFboII9k6vLrbCccPQFaxy17ADU
un7aZgKGcdObzxp2mTyaXxNLUmXiabiJxo54DAtz5jWIdtgPkkxawusTff7ZBTutY/UheIYTPE/0
PfXzy8XAEKeYsbCH1pt7RHHJFIK46Vt/hEtZwc3IBVTpQ+5dDv6OhgqBm4XeSBu/SuzjSBvifVvH
E4FbFYscC3wWhMrK3AkKN/YD3BN/WnYvyvJ58AW6b7jpDlnRdSclBL2rncUo8kUn/IBnRFROynv6
p3HlQ9UQcXQboPJX8YweDmt8vHjkK22Iaj8P1/y0TzVlXIqhYjjemoKMifQyDRyUH27/VBcatCoX
kciy3Htfdsa3Q849pIjc9nuog99slmQEd02O4gKi3d5LDIXay6CtHdn7UkcgJfhVsRQbjuC7x67m
61mvv90cI/7a+KqaxrypDVZpDyJzyQ2jYvnSgzwbA4YizD8J+XcSBhiwWmw87woF2IDvPe+FiyxL
kBKtUB/KJ+leHlx6SXVPgcN60D/HJF0NCLH1n+0HOZ6myhd34leW9T5IpfGCWOjbjGjcSlgrx/oU
QBLUf2ao3/TK9jDkl6lj8KOZD9MJNSeNRpbrrKZNBX7aZFNWIYTjbzdQNPeL7HzTJYuPV783cG4N
v1BCFbe7FsDbKndIdc3XoRMp/PWE9eVK4H5tn4nDOQdc0X3cDE4rxfSyedXecUS+UiciHwYg8x8x
Sk0kJqwKPFtTpsXUk3ujniJFIM0loz9rkQyOp9s3rkqH/UukJZeZUcouOtKkUMk8uuxulGJ/IVJI
lPfS0IMK/zbhWJB8xBSVJFxz7PmH0rsp4TL0feFAQUnCXEJGIMwxd1ATS6o6o0td218spBpraf49
4OUgJtjoIFcIB8ndSeKtzlpgm7eV9tBn3naGpMGL0fYiBRkxKvR/b4G6XhXY4bqBOHpi4KT6f1VO
yuAwd5XWpCD4+pX/uuVai8xlr/B3ZQ1jDiR0tschxSmoGHjACYZt4NWkeORJp0NNXGnPjg/AnZrm
OtOmeXRyB3EI2ghRqSxK8KwVD23y32wjVe0o0u2w2rMHIBsT5t+coj5SLu7c1Yt76qeSwDHZ0FEp
v7Wo/pmGXN8Wrvlm2kxOXhlrz6xv5DZi8vbC7ARB7CjA+OtBATgx14u5GVNF7Ii9jUY/oN0JnHcG
d0cD3fvJlMjp/gqd3+qpJVcnBoG4ukDi3Skn2pX+yM6zVf9WXX1XLWk8IIowB8tSNEK1UEapYfd9
iusBgdlZZGXZbdrIOUWfqm4vOJTeTmKo9FCEvHu5Bi479YQz4+MQNaeqV6dbVpDVUDBQcTBm5n7B
kduxIp3Xz2nzawZYEWYNmVOS9HxdVqgBop2rOhKz/WSN5N8q6E5etgsWpf8mb07bUMmuJHpoghHp
+zE7pmeYqJF5E2E6rbdS0pB5TtvUvRTgaeA2BltC+dhzZzuY7O/ZKXsKH4g4hPnSrFB+9ssgeez2
DDAGyeaItlTtXmEvXMpscC916J24XzH0dbdCQbNTCwmu1YaMGaqFiBvOeta2dUXrBDq7IXzFmRIG
MsmTQURhGtD1tZlNMmvSd/dYJZzGDSWdGuZEf65l4V7b2rf/pI0Ib05g0uREiDL3kgWogWouEbJ3
V66RVseIsM6PyyuNzsdhTkcHcCOMvtrlzU1SExNYdFqYhJgUe2aZCy5cKRnih+IVb3hWMzbMK/4u
o/YgnUDxN08C6vEwLOeZpKmpHXs3PL5rg4R0dfph601eMVfrHg+Qor5WmfXrMebMQBceBr/6DvDU
pBkPwWlKtoZfEc6lDuw24Gyi6oGJXJNW6pzNZX8/SwdrlJtE2v73pi6k1ZmCdOQxdGZWLtR3YQT4
EzrNdzjbSiemzt/lJTwDB7DJ3JtGe6CI5+ijmwGrXpVwRpNXT+Aq4EJ5k9t0fytcYYYLuqKjDXdf
Z6/hUphAr+RfaNoX0lF+5qGwIENKGNU216RqP936azqTZC7ByZ07y/IeGJBZgXVx8weWQbvJMN/f
D6QgoqI3w1zdHZiWv4LLJmDC/phONtzsBZtRKMPiZzf15o+p8nHvQ0MFArYzjrG5LuA0tyO5KrtE
FjMl/lov4pn2wR1PoJXbSQXhQmzY1gWGhV6rAyz+5oKnyuEquHv22QvVVYKhDz+tPPWbFgzWbuGd
SgBC4x8cdkwq/sWMLXT49gCML2NTQka5PFB2ep/j/zF0vRMcd+reE/KOt5euAP0DJ1bLor/A8Grt
kgzVAN+XZKze1sReVQ9IqOT8cupn0HtdVI6tckWJ9pxnPl8qMcuhH1iICzD+kGRvLo9UST6aGPI8
LeHiTiLEFeb0rdw33FVna9hqWlq2pb7fdkPILqJlELAAtn3YC5ASas30KkhRlGtOxVH7sO1Q2U0s
3UKbHaN7BTIr8gglVvmTlCJ2WK5GBruGhovMgJWEnknAL2ZuWWqxYjmJoCEC9QBHQ5lMiKEgVHJg
v2cjmZf6Mnt1SGPUpViQq2FFVbs79HguvjmjmlGEiZFxZ0XB18pZzkg1zETq6zZp+9qUMv7mU3Q9
cs7wM8p7Pr1ZK6a9eWEAHSd5g14bv34QAsDL4DRBa+3TCHAm20ifi0Ia4E5MbgzVfmXAW9CkNcsG
l3YB5GKC4oy273Z06JfWI8UMGiOgMK/MGFdV/Fmp9OQJ8U7LNOlnMGiWaCY4isJ4qA9RMG6/FY2F
E817eWm5/4LoNhjJPpauGgoc/cTpw/S1kEuIEvsVCHAQR7zK9uchbSnGBFqjVOIKp4AwrJupNCoe
XgZs8DFU9pataCocstdHC8326560Nw/WJ5HHfh21XMuKDBv5Xv9bdU9FCfLAd98KN5s0PuPbDHld
n5zmitIzinW88VAIyg2PxlQUIby4YgAalpc+h3xoXub9TnVH04ceSobGdYanSgV17MYfgjFdhedL
XrTnhB91HCyWKwkGig6QbCrPKMOO5BF2V67lyAKVYIOVCxQVqrIxNZ4UIAt/yJQ9WmoRPPDo2wux
iDqy2U0oWZ3GymYE4PT8UFfzU/dQfmN8lZ3xahFBZDsxi3N7IZUFy/wXnR/Odgqul40Mx965p8Ej
J7qH9MwXbAwMp31k8uZe7MJWeq0Pat/x9Jn9ExvBBGxysKr2A5jMt5P6yVi4tj7I2eji5oHka/rg
MLdnSD92V/18Qp5U9flxxzovvnA25Y5TvOWbI3JY8Osi8ez2oJ9v7CL9ajuSjDkCGSiXviQDyoaK
vnZYJ7mqxxpvcxBKjDvs1qIzy6c3rUTkHZQzMO6HHuQzThnzYIFyrkFhmGq/k9MGWFh6F1B7Xs2m
stoCHICTUxFswbmd+RBtZSB5ocn0qO/GDi2d1F5XiKYVgVXo8kFmTekRYN61ahCv7YISeaEZvhkr
T9GaM7DM0CSbMPt4G0DX47aW1hFuRQ/hVP59k9ClfL4Esjed33AXcoEHB3CyW40jBJTXFmI6Ppvj
w2EmFY4Vmf3v4YR+C9+PjtzbCi7A50iTZDT9BR0d4jYOApg2XSjYo/fcZseLTqGCqcay1HxnrOoN
guS32R4NyamveM/e0NTIg1xHRpbxJ+Vn/0WaX+hk2NCs7NdpI6BxoD+Pl9CV55RYfRYK0R65UPFM
Cwy1OIP8Mf3YvQZjqb2DqDhJDLRvIi64Xr5wWxgtr/OUE7oNARRj5jmZHSoQ1cBPYam0C9OMQzlC
lIkAQ9PH7NpFBD3ceXXFAyIwNlv0kqv79W1DMwKEoIpdCQTZZJuIF3y9L21XvhUZEt/1nVor1NzJ
Ecn67fL9jWfbsK/VcWOWWZnhCn6rUwhl4swj2ImueVrFCEmVLb9C5I0yGGZlEbPmYE1+vcXWJlYS
EPrcyZN2Vz+ilSkeK736kohMrp6/fAl/2VDU9tTJ54x5JrQd236gqufAz/zn6nkxRmPGy3DOqjUx
vzGk3cOf54v45kPjW4FT+of2bdUT3ztRtRqs8Ms/Mmf/I4Q03IX8U6RGF526tucSaGVHNYnsBo6X
1V1jO2W+0Jf1EoNQyBy+HMZBotw2RgDPuVjqQ4590aqWi1fWZC25Qx9SU9H+3oSEffZ0hqiPqp99
bGORHd2cF09oc6l72e48d5JJOrOpd3SK3pjKO6Yvt51emxegr3/4k9lD8Se+eDQp5uc6IRiu4kt5
ZRCugmD3eWBWZhqbVeDnbFAxN5zfn8HyuxnaA1NCjOdjbMvdAUpldY6K2A7wgjuziZNmi4WjC+bY
ynhF/1wk9GqLPq4E2Bde4uc2pDeYqELRKkYzREJAqjBRoHzBO9feDBSbgGn7DEJqEzLFCz7OdgUT
+Ul1qUO0HB4EZ9vy5zH3VNwsCQg81LMCyk1uPPt8dEthPQmnyhZeNjRi9gxZRdmiu5H1Fy4fZTtL
S1BRcXBq3QUhHISDVBPhRiYOeOe/wQ3x2qTrGMHdwmg4EsQL/P2EX12RmB8/o9+/qGpX98mcVccg
rWVSRFEBPFHhwCZWKsLjvHqvGOhglB67TIj2ldYKqdBO/m+fNdZiYyN9VXuZoY3iNc+hzl572pfX
26f6ytZ46YKu93mkwCc8J4wWxu3AkX2wyLh4kfieOovJ4jCH3FUjVb2CjW5ECE+J7aPVAuprjg4i
BWyUUOIBh1pLLAP2Vhw0zXwb9QqR+lkVSenz0AkDBnfakl24rjBGUhRh8PQSATatcipAvK3+Kx2A
M+HJi2ZgmY/p2dTZ3TESs56ttuLyOUqk7h6hGy9xaozXmvHVBvX0FOH3YB0PKp0AUDQZ250z8+mb
TwssO/Ctbk6Q1fQ/ZSWWOXtaUYIlNgsreDxbrcS1enW7NA1H0SOx2vV//CeJB1LUADTymHS4V15t
oT9iD0WR4ofTVQBMQ/YoXFfHZDwZLStQU+JaoMrEfqHCpN3XCxpSjGeYMfIdzYtqaMeObPXt8fEl
vuPDxTLpBUxdhIQJlNZj20o/ybAmcAyv96dJDjW0eThYyG41Xa3mhIGHn+839jrCOsGLSFgxlSya
7cepiKSi01Yr2lfRRiYNaYStahZnye17jkrWQncCIPY3EpVUh4OJ3uHxWqiwCqHS+Q55umkbwph8
dZ+HLafvU5c/FWxS5uqMAyGRcoCTpZb30PQeKE3yV+X2XCZ4ZvAHJPsVGfUdyU+NvEu0cneOxMfl
RSVFa8Aj+xJhi7DTZv20rwSHFFOxhaY/IS8Y9KOWi73k2kQB7V8RrvY/BuAmvTmAsIhdgdCpFF4u
JyTSg+qWYo7tgNUZG7kUmypWkfzxibhDKvJ0wrrW7Qg90txtOMmfNAcGcInHX47hlcTMQN7kcrhe
thWkecded8RR6np9RKUTAbhYiNp/lbB6APNVi/gmYLeNoLX4r++dkoXs62TEOW4PH+nPutbux2P5
6cF6WjjUoB2nUe4sto4utp1q6N72Yq9Q+mzis5cWfS8yhxKiFK5rxgHMAP2TM3ToquyGhqrZ6mn3
U556SjC7soCD0yhsGuNHJEMbRUFveuDHWlsV3GPlxex4hDwsOWQCkX8xEdHqQK19RKzuFohU22J3
vaeFi5tWy5Izvf4wEN9mx9wSew7kcDZx9mGvvAXC50GAwQ13dm7WMki0ssz1A0aEGOmkG7NhjF81
0f1FmZ81ODhlAOKScuEkmgSKr4RIAI6CebXDkLhtI0TEo6BHa48SSkvlw8tz97mx6KvAykLsRsCe
kuBLSwrUsUCdcP1qcjIs8cNNyM6gAfQcBCFVmXLA6cfRUOOkElsc46wLvQ3GXa81BVX90ZOwo0rx
S4eQz1E80EsVC0S28FL6RKp/HUaDoOLq2lLxgNdlLDS13VjmHYJNXs9hvN7L15/YdgmSfXRTf6OA
aveuhqOaLemVa4xQvgXiRnYe/pQ5FpKpbjORukwqaihQBg9AJDfnakvGiBTKLUX3wLAK/0b5BwTy
NBceO7viiK+gMUwhEFWhA5Z+zxssAMh5H8JMaIPoqdIwhS+OUvbd4rgk5GqYg/FUdJPK5ML05i/I
b05MHAym1ndyY8+dkr3OeSnnItzyXGaI5UTCM4njTDtu+yM9/NjWanMEH6OfjY+V9nTw54JYU4Kn
JF4xUmc3dogo/wsQqloumzAhZ77aUpAHd/juwu7DGPQCGIENgI3R+C2y4iTyt/P9wtjXYef/WxmV
21jmoIjgJDFeDZZ4qRO6t+E/ltUm1WOITa9Qnv7tDGPR3zu55m8WMwha5VZTgiJ/1IPeG6FpmDTr
O7Nb802n4mgnbQaW3Mxf3jmVmVMUyzfnAvSIrgAyzajNfar8/rYDWpLEcrrjR/MEapYm0RT/MuNv
Pwaodmbqmdp6gho2zhvL5KZzhrDVSGUiMQ+z4hAk78zcQaALxygAFXXINBmGNGAYPUcL8dSZvmNm
exnQRdmDzM3WbhHDiikpxN29HvNH2Hrj/Pg5IgAcCD4JbPnThcqdhZTEbDUjUkZ/jnkhU2LfkiPJ
4aPD47nbiXSxk2kI7+FmDsVy5h+4iwtmRiYHfFPTRsj/Td2HzInfxKE7WavK/GNrorugRsdKj0S8
LpKGyaHgxEckNnjDysfm+ecQ0N/9yXlSnTkzCpmZUVnX3wnqJPJwp08Qtu0haqIBwmiZBxcUKSrX
9F7zokh9d06G3ntJgKzvbeBADRq3ANA/EIR8z8bAaqb7yDiv74ewSLISJ/yBT9nCUJP2sA4yX/d4
qFQPFkTjc6XcB/zXf+Jcq8666pZllTl3i47uREAiQbX0aRGrVehJUwNpbkkz8MvjGW3EeNqlgupG
YwuW08pII8eSiobXP+Uc3OwJP0w1bh807KFeBVLSi2t6KBz4OhIzJy7OR/3XBm8od5zx/opkoZOw
IG4nYfDvY2+ESFXOwk6YhjaIapTjIZ8as9ggYKdCpkmP+TCHMUCoLrKc5vdu15tCYSYmLG7tvBd0
oWtn80RFXcn3DDCzpzJZDNNOfRCt9on4EmKku3vdmnCyOvBKqUsL5wBA8W63nfWzbu/EKmly3U6l
v9qktH+z2KwDFN9xUZRwpmX6O3P7G0n7GW5UG+qAk5iDsVDW5OuR/YjEu4JJXrp4Q1i3/Ze7qwDI
Az8E1Af+nmojG2/oTNHskKdDPSs4REvJ4LSRyTIzqfg9THP6KA+OPACC5CLy+lj/ADVcYbQAqtt4
6oKjOQ64mUK0lpMF7s1VR0AgoNsuPC3OG6Fzpt5Fp8JeKvNNbjKIQpSPFU3cr0x2ApHJ81J3znWT
lP0xqpP670+60ncUX2cnKyASjQmJCsW8QqqRMmJ8W4jYD5L6Fd1Bqg0hzAEIlJMEG/aFXW4Glly+
nUOjaFY+yWbLPFAJiHzOygDtOIhxudsu3EZ4kRqoY9Fv5nbcGeD4JJFSDR+zt4rFVxEZb7YyjV/4
f/Ukd0bPNuCt2ayfDrTsNh8vZlKcfT+HnGr0tcD9odjMStMbaurO/YTVkWLtro1rg8eLpGFEmdiK
I3nK0srAPKJ9X8mpOdMvprZ7L4Oo6uC8mrxofd2M4l0Li1B06Tv2YmKZ7fosU7ViqwASdzl4eko/
Q+iw2De+P3ybdKo9WyixEz94W6SiLZlMiKiAbH+U8kbeMVgozBDYFh8i+ttIFHQYFES9gNv1Qc4x
2wvDWavQbw36gRo+PstpiY7yPjMw5YXjfG5zyTXb/jtcrD3YGzZvJRsQpa3o/3cVbJcsBd8pfWT/
kDUHQywezgBxld2kkdjBv7jkYhg+8ZbqJCEPc8TnTCX+I2grmcfqkr3pg1bP+VmHCpNpEuV+B2XA
anZ0Rb2Qn9xHwahJ5wmxT+fS5//+73EANUJtJhOrcFse12dH0kyeXRvl0LKcDGyWITvjc4lF0wAD
jT/UWoJqyMlVRhlt3i7XSQiH4KPjVgrjk+8jO8CL2AP12xIEkB56HBnTI9qqQDc21uoD2r+BuEtE
CL+P2xWTHzAXaJYOvrrnaeGAhSWVEueDmuWRY6LCAHGUv/HbNQ0LgsPaabZGS2Vnb+GSOvgcP6SJ
yEHFB9uBvzhMck3gQXucsLWsIqQ650XgveHfieGMWIdGT62i9ffhb1B3GJiyImSHe5yVvgmWocwa
+ORb8tysHD3I8rEtxZeAMZYBXBSvol3tpqha0nownH80mDQjF01fmfx8zWjU5h3Q6HS65CyB8Zy8
l1SCXQyQQ3jYDyfyFYctAZjHOssZbOUCTbIqLpoCH3FMQQtNhdxVU8O1XRL1mqHySmkpv8woBWxl
0J6RlE0+XeQiZDSQuzM89Urx0rrah9GGQwd1xOGDh1vNF2Z25romtJheMBaGiJGnQrQ8wJwO4W/c
rfI61Z09/SODLj7WdaFuvo8IAvpaNNfQ+lVBEXf7t+4EMQ+Sfq9ZrF5y2W3BAN5xQoB7EIqM62Ia
I+0tWVqN3fRqrfk+76FR/kjew6uvpssrCuJxz83/5HEvnvmOpPlDtoj0lrs8smb35tmo3AHeikUy
E+bkTJvIVSbB3xYimwe1b/qJnpx36XqB75q5YvDok4+HwbjR3u777whTsa83ljc8EiIllzYP6O/3
tpLMvZ7p0BwwCZl5aIi0xIZAFYWm08jq7g77bnqy8RM5hCNhpr2hoMAfN8cDXNROmKL8xmH9rots
kbtmsvCEJPNGNccC4mm2XcBwTnyQ2uGF9gysUqce3IWmqpujI4rwKTpHRRMIb3PPkmyI1zTCtSDL
AZXNEAKWbAiyzF2LBX8T+IM1RJTWz9LgR8monoui4wgxpG7G6/DDO2PsPLUggBGUVy/814/E2xJB
Ftjk3vx6gH50tyuBjxuhUv6QPrGdp4WyOA1YZsSihQng4FpY/sjVYIuhEtjsSTnT0YgY6Fj3RugE
3sYZK9L/NjVcLVpvdOFWz+jfhR5eEPk/2r95S4r0TIO/f7J66p3opjcN3X9oyxsswCKoPSAN4d8E
0sECoPYAxeXqfPzH+J8dirKmy7ftATgnat4iwzDmORC+9Qj06lnEURVXhT+ghUlMjwMYDHbHSEMD
PBM9VWZqRfruNs//OBX7MxjuA93iHDZqzxHerFL7V6YoJimYwWCh2EEv6aUh/pysuqKfYS0M8fJ6
b9A2JXLfK8rz/Y+73aIuJVBrBFFTMmvuW1O4+FJR0QTjkMyhs3l8jQMeYWrND7pfWgJUXufMHpYM
oqiFbwfDBaFP+X6v6LpBk15rfaDa5gAmTIKBOK3FSeRRF1IqhTzwvEczgUM2wMobL1vsby6T1x1M
+Zggd/rXvO2raOEZZ0extWiwQ01kCoRfrd7sOwZ9S+VvcbiLDWqXCh3SoVKUag5fDCe+IYpNkGcq
ulHTvEmov5owZTxOpKcIz4ixVJsbFVDh+u2CDDuJf4AmxHitznlsyx6nUz1IZYV4oCMm5AulIcej
uou79s560tRkKKIgvXr+kmLEyvZjqrJ9EpoQfw+w70cro3v33lBxWP6IPYX4CK0q4CP15yiQIrf1
omzwdMRaGNfhgw/jW/dcxo0y36LwtGXfF41eQiOAWv7XSMXF80Z8bj5WwI9OMrWB6Zj4I1ECcti1
U2kOf4ya1VHMtW4MvJK6bdCF616pxICmkIH8m/DttifBReoD/QDOq4tkM2QYk91YNu2BKK01s7Mq
YLFeONKyZEN9H4QMM6y+wd00fU+JXxl+y+DVvZkHmJH9arLPco/wIhEfrTj6fjlpSVCuPAVZtVkg
5tocFMXd8E4jMyDZE7BKxLVe5z4uid1SADzmDS9riLMUMH61bXLXVXDLoKU72ygZZ8Mym3GPhpdT
HSMn/gIDkr5FlnnKB76y0+8OEoX5cliwXI8saQWuESen49FlxVvjJuHuHkBbDYAEKVhRU1W5htDZ
wa/inJ/QWzJ5CB1ie0xoePpZP2Sa2dz/yndewT2+pWW+KihU++2CcTHJJg3Oj+UcoK3IYc3KxUg7
Qf3Eyd5HbpA+ZQNdMK620awpSWdvfsp45BOB0Dvz2zTEwthM5gPvYjuR93K+woJD81YeydJ8uxtv
J/nRAOPPZu/OJ53QV/e/LgZiURxDbIoFNQdhrgUyNqDrvBSz91zDdh8+nV6zBfG7LAREHzsYETMo
qyj9cf/7okNrb7T4jpJhjMefjNTylEnXBalRCvqQZZsG4FDoAfvtQVRGABniqNW3lTiJjqSWp5bk
bKfphroYTEbwG4xqVytVMGIew/zKlSQjHOh4f7KG0vfvU2w/ShsvgXTDrCwEl2fQG/YRoA7mWIXn
XTe8yYN6mAR4FpSpo5ex92sZkvwm+UprKC4/NMivC7RDnHHt7EaW5b0qSODG+ihzuYIDC2iubXay
/6C4gVjPSWh5egybccUw3h9HfAkE08BaFugLlmn7lnTk096nrBv+94qu3Y2vnucb/3Na7AtfITgO
Qh1ya6f3fahIGOn9Gn0147V4MnQ4juV5FSfy+1Tz+wct+gUJx17kU15aaqTQuL0ydf6CYiymxN2e
LEvAqMRYXJLyBf37NB4s/0alQFJ5CddM5cdQx/JPO14WgT+LJAMat9IZKvP8QXsBjH2aZMCn/b7l
87Cqr4ed8SgrJwZbiE20zQAykYBAXr/YV4wHbKnbcBFbziAG+QIj4nlZbqW00jsT+KlGaIg/LQQ0
Fh6wsfhx3gtuERdge3qU2stvEDsYVw0C0sOl9ij2laK0wuzUX01n3v8x1zDNZHcUOcLuUx4+D3mJ
3bsWWy/fzJex4TNYYDLrZwg2ikaYQLYUFigfJRXNJBbM93l2C7OtpfSo7DoY0939zZD5vVJ97BiP
OADPtP2pQ7dqJyX9d8N8ZWyi6ChWx4tVNp6X/MWjFGlf4c7yZaOCiovOl7dqHl4WKqCfU9x/QR9G
IJR02PMUnHHfIk1HjjLthl3bh5+zSUZ0KoY3Y73REdWi6rOEXOPZ3ZjhVPo6vcj+adgWVCJ5tcPd
7+tj0QHvClKXqbXvgbpiIM5en8O7MhqVmL0MNkGn+OLcHuuJrqxSeokLOE8z39jm7eycz/QFbcug
CTUwGVJux8hFHZ+aNAJIhvY5gMu18zG1/inv7tze3uw2reMCCTkBpSX60NqqDE7u5fy5JGzptYbb
gWzZXjyAxrRczXmqH4CXHAiZmLGMvT8G7xHLj9Wy1PMUv/ecl8BHIQTk8WRt9Zam2MiShyuU0Xjr
r91CxCxRdyi6wB4vHJO2X0xqY0s66kd3VOAii2/keL73Du/6glozxwSk88UuHXNXyqyTdZrczNCI
K6OAVtimzXP9UtUUCfX3Jrir8pasgLRRdbMFCuPbczMXmkXkJGB9JsIjDcJmyQv79KmDNMNvpnPU
uzGGwzpcMOgssxCMBEPjhEniWU7OH5visggNxeoUMXQSMWAcFa7fXxMdvuAT+8kwzbt3H615kX/j
Kbqi95OPMvhJR3vrOY8XuVoPBCAw8nSH7an39L6G6UJ0DaOvJf7uaE3h4rgbDyZ5cL46lG6WwcCR
8NJExEj+fErMXOwpf+VGPqeeoqWY37o5xz99NFp3QYUAF433qPsGvHug1wA49BsVA64RnOE+tRyn
hM8nkfhW3iFEcDr1voVC0t0Th8YLmIu196L/Kad4Tiwh3U3UuE6t9qEO7wSNJXwdqRO5U8Ksds9Q
abcRbQmahsAzQq30rnyKpORgftD3AcpOUJouaN6O2lLfStWQatIKmOujj4eC0NBgh0XKexMUSQGD
yaYKLCZ/e0fOK28iVZCcA0AzQymMm7OE4Ep/07x9c5xr3uScVyRKw4vpzpeKKDA+aD395docd+xa
HJs9ZLKtWgd2Zb5EJgeAKanMoHsbNUgaSP593gYeDaXPR/au8nhzf4XiXdfe6Wgzm4hM09BEMiDi
yhuGHQeYhJ8j1FxI8NuR/FKCjXLsmX9XS/3b7ZWGSujnmxivdUkeBBebmlJb/za9vBTtUly40r09
TLyzjPyHfvTr/VRCmD750WSzTqAt+DGkF/drNbIII2oPDguCz3yHbGYMXAUco3bdWIeuJkyg+N21
W3PpO23irvrLWgHiIU29WQCkOOX1kXGqE2uC8B2F8rBcJ7dnCVDovmJab1mJzT3hf8wh6vv9dnl7
zuARcQajFFHrZhNXvDktcfKWRbkdWxSvJcQz+oklMXOroUcoOEMlRPptrjnWAbiqK5PZWtENJduq
dqwFJDsOhaNIEkb9HpnfELMMushhM7hfskA3B7zaviK68z1zZWAzVuOvdhkSmf6qp6u6XPVb5mlZ
XkSWLzj6KU+B1ntsB+OIyiKNnNCArEBMgGim/ChMyZ8Zh2BXks+CR8orjPae8XI/OqlngUM2sCCh
tSmgQSPizAbhzlg+nCUA5+MYc3DuoFjyybiviGCsn3PmVIPk4KHy9v29y8lj00bz63sqJPJU6yIP
ktAQlEmvf2IHFFXMeF/E1Ls56NtkU7i4V6kHTg9++u8mvw4D2O+SGOw3AhqkO3eVqvs1Skb+afLp
asQod21R4CaL8TE/44FNusWeWGp6wu2aCHBstHB0OX1jKr3rZps8k3lVgZ3bHDonjPdr125lP9Sy
pWdTteA3XwPgWzKCJYGDU2zjvTjsL2GYXwyrEC8Gj4iz/iOtQop2/WZjKNlBvzFLYLPjMVRdoEX5
2mwUXpOvV7I+tpicEk4n3xpBAIHt3tsbQZ0Yynoo0sdcqZBECxb1KDtXTlRWJeMQwglnLkR2rmfS
StugdQhTy2toU53V6Ncodeqjk4ynkGMv4zP526Osxvge/ASS+i6K70NZ+IbXre+jks+jHnkTfyJf
rp+rBeN5NUIzNuBG5jjGoi9CTgjBbaAY7Jow8XX1DZBWzgIWWlEJnJtplvCDrEutgQFlGUvfRswq
nPTsJJJ2hYVPjx6AVJJhURoEtkCrteStqRPXKqGptQNgXAalJvtTuak2GuHlHN3DP0ooKDXUqKl3
T8VXK0gGt9FWuqhng+4fClih7BkW7fhhlCg9vZeR9LpuJKHPt5oGdf3M3JrZDNIxc3vn49yyd27W
8L5dcH81RYSoRbt3d6Js77yHjzv8+9CXWgLlYmjNyZVh1mrmaq9Cd24nhMzCTcMqfYDdt54fNm8D
Fg8n7mDXT04UI3aCS9pwITADP9w2Vug51bygb3ZhkSmXpAyjW8hQXFtfrlyu4/THa5mNlXVHF4uB
+9GFr/uST1EHsZk3pPN3RSOPm/O0aCND6A7TbCDn3om3p6i9VyrrvQhkh/7cRRrUC9mAhnFQuEXr
Ldkjad53eNHCRBnrsm5EcTDX8Kcm0TftkPvpruMxw2rNwxhOadP3qJb8Fu29dEKJ1BtLqNfsXDEw
Vmc52F5qY/VOJsA0AW+UfF6P3aczb3mmqht3l06J+VCvJh/Xf11jNXmZLRbOAeQwbRc1CsJxjWL8
2QLAw9iagFDy+QGa5+MNNdoqzKBiTwHhAUdKGOIMXo/mG4KTT4FotFopUlsAtNhKvkkkyiGpgYc3
epWki3nmFeKaQkFogyugS//S1Msz2+9q2gO0OpSDHX1j/FqXHTk1vLMqK6EGqb14vgQAcUxNzabS
qxFxXdlszA3GljfoygLMZDI8tOkXa7+Zi9Z+e3Jz4vH33hx6VxdoUNtu50qRNLIokV2AVADKddar
2AUgRZhDF88dhyWvURwBWZk8REODnZifXCFcWteJ3lS3QDN7BaD0Z7SPCh5/YQ27upW4QqVBUO4M
al+Hk48uWwTmSVdKy3SBvK6+ZZ5zy510ymWbmc9mO2l92H5SUEJBJ21PhjBr+9vk7eCoTRBz9ZYS
VQuY9JfN36DPdZW5VCr5IS+2ysDTIwPIs/vJKzrBp8UGUbBtKDu5mkHyyGdLeZTib5owEdemJrT6
7EBXMLNNy7M/dB10vRN8ckfkyr4wVwjVBAy99yqWus2tXWPzDaZfMqdubQoY8d4rjQtYHNOY5pt7
aOiIQxgbatYCncI9S2VRcymHgaU0Ziqkg6lnHBbUC9KGc+Pm1AzHOVeVDaT1FsdWjDocvsTXpELu
e9WWRtzavSuNJKEOw9I8rb6K+WIb7uyZT0+ZbzSscewstZZ2SGXYK0YmbnMj8sedVuOJZ+C7+F2O
h2ZHvYOVhAWdwB5ngltlmGoVW2utEEEQLkcDeN+FTZ+kLKvjLIb02LlznGkj/GxcxpWKrw572tMT
3B/Q7akgb+G8DJS1pHotxnI2XDctwwsYWQDnk9V+cS9JwscuuMZ2Of+lLba2UH0qhBQnVL8eEnA0
c2sxv5XrVcMC8j32yh6X7o6RUPPKui+xHaUchkF9xqqMcAwoa9W8FU2ahkcJ5sd28ac79k0PE+L0
LbbYmlWz4t/9CAeyuApHLbykVzT62wOEsDTSVEEhRCp/VJPZZCSioxQ6W8Hual2Rwx94DuIjNvuE
u1UL/uI0mvnY5CFZNsmXEyjg0b/uo8KmQR1iSqK5+1e6vtXh93J2f8s4AMbO9WHlnOO5svsP5W5+
YFfHB4tsujqQr4qV1cZsVuUkDGnKBaol34OKyRNCRQ0OVYKYbm7Ze9hpED8/suiMx76qzl8uV2F9
LrjmVQfyWLnDUdSt04XmQdiv/3sTt5U2ztE1SFpg0RSUNTt/NMzUuZ7G1Q/dTye2YgEOzq6mYkbQ
q68RVn7hCVDlhVe4zv2xD1r8CPnl9zfk8fv0pZADe7UGD7uYa3gxfydQA6buywX/irdVuUqqTQ7W
fYNJiaoFyP8TQfmyLACaodlk19dVfRu975AvW+DHctyMqsLnyLWZVoIXlpXfB4vER+HkiVycu4tO
VSe/6C2LdQhyHUdwjk4kpFh5qg/I67c0BGoz6n6J6OAYBOj7+ZEdc4DNKnRME50D+GpCYMSJWs/e
60cWQKXvqO0aYVMgUNbxcJ1h9iJSxGandJoyckjndac658uyq4gWx08cSVGhhahWWaC2a7lyC9vS
pKBSA5vWMOupL2G1bkm9Y6didHC/PVL/JXaScrZJs4t3Gn5auC2ZvY2pQp08Ptqya4d01GAjyzCQ
lIQyyck52wPAM86WVGwgblwhGZ+DpO+XiN1/0PofTEoDcFyHavjJ+BXrgvWnDNO3WCFxRFRhNy7d
RPO++3hHRsXwpLaKPdIB2uYqO108QV4nLGkTQRYiWzyhn6PIz/FxKGrVi+dZYgIM2D6jPbeBQL7A
g/dUWj5atD/+RzxKnBSBPfTASdwQCBUStiIw8akxmn3TEE64mASu2UsAwPSintvSeUfheHvJ1B1u
QQG8w161BFlRaMCUIJGnrHnzb+JX+f9Eb3SzBs6VKjmRWbnRPiTYSpv+x/lS0CGzEx6QOElJDG3S
38i1t8xcDdefxru9yD0iMF7dzCYINUP7swXNuIMb6d8/dnsA/GpirUbh4ApgdP7pKzXsq4W/J9gl
aVAPLTUXDzRLUyg33qxHUkKyweNoLbK5Nr1l1ZG214Qkz+3NCfbbIqi4/B96DnaKue5kF9qmdIyy
9qrta8qOcTPvQS2/Cwagz6pASMudI0NfZW6hxa2i9e3FfSeJdStFTnHrYu1/Ja9q7GO+M1y0fetH
kG4zCNjUTHJKEYSyNG5jUrcEjKuT5S7npg7o0CYjepHP9LLxlx0h8ntCrz6hlEKyKLsRO9L0jW98
kx8tce/IG092sozUylgaWLVBW9e2s35gSRTiuqsp36y8EyaKHvW8ECJImjq0yff2MqpwoqEB1l+P
H7GOK78L3ag8pSfS4KtqgDM3ucmhXmGN0OyYIziI+/FXEGGNkUU6n1LvksAaY+du26SMfUo714e3
4eriI3ZS8TewGHPCijmt3u52b2KsUYtNLmvGxwmuOrd3garha7XryTkH2lzpx3FGekRcaUsYWx9Z
UxIe4MUTuk5pOcOCWZ+dPBp339+kTBG6DZxhcpVQ+fopOcvmdPkoYb5njdrLtowkaimATJMWC3Jp
YtJ9t/rJD8/RExKHLWEb2n5fFkcahp33DyP/+hLCeEH2spbPS2hijnhcfoz7KYolsoOaDG3kQOlN
QvKJllSgM0OgvcMGwRSgOqqAJZesgMRxDt5Xj6PXLvkNOR8Brg7P75aQPdN/5IhaN4jncCo3lIzZ
X9Ql80BBIGBauWh+1wv8pNFkt/phetdaFvZ6Gz4FpsBMPxY2wzHIERWM0+EMEaCFi9yrhcjmMa1x
GKf9F+RSz3RapYlippQg+e4yd2TqqHa4lfXg4wt6TChNDmUUZ6vKmzPufBi7y9+Rt7HPezeH1Pyi
DDJSW+h0G0dH4l3PAHimRrOqhl0Qun5rtdzSdHsjIfvLsrImet+KX3jLZ8bRGsIGW5ad/TqC7r1F
XcteAsSt3+W2SyMoyBJOgtzPKRYZFLwQsi+9/0OrQmUL/aZV5JSHmfc52dfZryQCjEmxGqi5qCj1
Uj276QTlQKhoCITZcVqzumRb+rEiSVLKrit9pjcpKJXG/o9l8M0NW8YVBGRf+72v/oBYibxsTDn2
quGn1IdVDvX2lfXHCTW/u1qhpAS1A4yxaNiUc23vTQk5r96hGRTgTtj5b4CkEZD+FtASs+y7YoVA
aA7AYWoWO34Lg3uS+dqBfaZ+So0rrTA9vjX13KHGlH5Cn2FYTINP493HZBJtm68uIoQma+zIbIo0
kfRWC2TJ3cmIV3LLy5CslHzwzAc5KEZZ1ow7cFBNMYv2gmR82fJLNqOm04epHQwkypVyd6F9qn9r
vlLxeHpzRhOMWOjohnrU5p7xPBRDkFGcoTrsxp1loHmgHAghL+aCHx5dKiq6JJU1glaMYW7PbxPg
h3iRKNMexOQ2+GihtJHutXQQ2zfM2bJoG1H4SudSErRlQ103c5JrbeTtPxsohaqbyh3dJ5d+f+wK
ok4022DRAN6gGpSJeKtY5YqJNnbRkfkRQzVbxlg20L+j2PF5A8tnmTIz2OESAyya5xh3uhmtxfG3
26Pb/2+jBp36A/EOKQdy6ommGNdrCPvXhgHUp1+P4kE1AZDoCCwZG4vDhL0TERHParzxOo9uHBhg
tEBmDEfZWT1J7EkEbFxE5aX+hxfiayHmBEPh5xJzDC8uhtpUzrOteeA14kKEh7GzL9hTVRqX3kTr
XXuatA0YBlsvgbn8oQCs3swYHkz8MYJRVnNo8v1ysumEhvKXdlffI96qdqk9kBqucPh7Lpgwl0Bd
kQoZKef7vgIylh9DoAdaJa58ZPFuipb9RphjznKACc5PcRBSBJOj+tLWILSbjmOlBh4IG04/rGw5
0o7OcpUlQju6VPKIbe11DWE5M0w5naba3k0PcsoZtNWtUaMn3uE5weZUj8VT5wQyxDEeoHjvBssu
Kc5E2yoVcACMfecKIb29ZH9B6mEX4oDGXGtKhJwgWPpr/Pv2yGARj8v5UVoX/FExEEZYFGqTVbUK
EAnm37Y/2tym27keMLn/xoiJbg+Is/pVioIpujYd1OPUO5GQqEO8q6jRyG4219ExMsfra6Ur0gtN
ZxshGmrfFOjhhKuQN7umBQTaOpdRw5ayQ6nLoGuvsaY9kpCZUHQBEd69R6LJkluva4uRjvY4a1ph
RtOCOmGDmF8+KBHgf6DdcIlg4G73SdrEaJiBzLAu1D7oSOh+gsXHzqdo4JLlM3ZBpRRUuW6iCiJM
IedsiEO0wFwtihCvjvVabxaHzO5D/i9LTPMBnBhDvIaY90FsYSj9hdRwEzPDgUx/BWi+6GwI+oIt
PfjzjQ1bwjY8nobtguzKE40QiAXhBZzdGO8Dpja4qImkSD8i+XsAEv5eoitQEX40x6e3vKw0KjSW
JMB8jE1Ofkg7YjWXqoDs6nKW4xovMxz2yQyP4P2w1JEcnyUJnpaGc1XlGNWMftIAZsCvV0zdKtzG
E+Z5FE7zkHvVthuwlij99HGSt6Ph0B+d9lagWIiAzPTJXIcXpPmz3hHxAkPZcQQd12EyO19YT9gQ
4w05IrN9pfBS3XUdIbZDw7rEy1bM834EOXHEs2D9nN0bCJaS5Phpg1O+rYVbhi6WZ9RN9RRsZvn0
9nPFIvi6Wd8AxoCLZWaeoIE6HJ4glABG4+a4/xNnvn21dTNWfyuQGk62s/2N3a2aveZGERwfh2M3
pucOaUhISVxrhYQlGNJycNF1yWnokJhjXome4A2+ULFkQ7GzMNFSl6mHSvssqK2WAgXRFdg5sO0s
XRVlqoEKUdXa8SVIMfel3n1sRFr+tYtjwXxtG0kOlNI4J8yiwFbKkNkPwnf8L2ihWmxaczeGEJV/
xHVj5UNIasnv1AKMAZtScGk8UeRgNnvB9RQnxvGY3ZIxfXUZaq9pdqhA7xMUNqDoMFxOQKm++sgF
rie87tcciaPnaIFGkgUu54etWm+cMuhZxNdrNQQnSNYM7DM4FEzn9vLBWYc3u5zqUMMvbvzu83z+
UhpS6GB18VJZ8SQkNomvm3fsmAWRE6IXlcgDXQsqDdTIuOLfp4HCgmP9O8AGKj8QBvf+NNQLIlbX
BGpdGbX+64GGaCQG5k8uSl2hsillVFMTWErdvZ5AZC11fqR1Wyg9w1q+bpU4tt442hRhwew9jafO
YJxiR9VIfywhXeRefrmJDo5jnPPJcGIBcPedE2+9D/LtdBhJByGSSCyBFspro7XAbaGBxAmZXdfR
cxcZF1SzwQG6X/FM8sobPMh6t4b/wImdn2djXTSswGfG+MCBA9bDVjZlZJJwXAQgP8m6xXUFe1N+
6z929KoLzoDR6+Me6mQyZMKioPd+zJPoRdYsN4ylX6NCGwXSoW81iad1cRZlDDYAgioUO72qSqHT
EFgvIwK8tsSK1jasuOuFwud+gZqu45EesZiBxAHbi/X4PkUAxmzpnBB2qZOVpoAM2zHLPyGSSu86
9ZSCiQjIWDNvTEFctnk8WI5gD79XgKt7n07kVy8STvRbqjXsjZdQQPWr+Y4tWdsonchPWcV1fri4
wP/jC3l+66rEfj8+X6Gdbm0aPJwS5bjAGOt8BFf593mzYMdEm/4ElGutBtZ88B4MQu00CTnB1noa
UhI+2OUY8iuLkNhOuGpjaagfLBQXea/D5dN7gEobM18LE/7fZCnPIIyw+P+GnJYtMN2LjAy1qxfw
fP0wt4cGLCMI0Q2jveZEl7/6AWvcRjr/Q/miYQ7dcD+hzA1SBA44ttL/gmpcxqZLUTjzQEcRrT1F
dfSffb0eIG93U1POot7BUCUU5HeXlmDN4D9C4+lDEXQAC34S/vTeZ9dLdsaoBiVJEuYYyZVup89U
7Cx6pwaL5ScaW0Saz+MnZ3gb3AZnTCoEsgbvCu6W655epqCPP4r0z1arjioe0a0u5vk4z7e4zw/s
AvcwSxXobPBhIsbBCQQx69CJQmwsV/nH1Cn2MRa2aywfqR7rKPWCSuRREPjbWPQEw2oXzElOiw5l
j4yvw+9k6vin2CLKhFe4XkfSx+zJF+HKgGgZQGS5OsvQPa2xVZpFtfLwGelANw7az2L84yW8uK8z
zQxLTdloyPsqK0rZS0z65KCjg+c1qeVXm4h1e8tV4250Xk0uGggTrKq6LXHZYR3B7ZFCCBxNdXJT
TvuioFbY9s8FgbEJ0zdhf9UkaUY1nVIuZf8lnHEKYGwIT5w3flZotj2RmMu8i4LFLkNlKsq2Chn9
BQMtq78lSUe5fbZZbh0AUPxm0g+dB3KXNTO30Pplg6RVqSn5VJxC8c55/IwrOhBn4ejd7vP884Ab
p8JIV36pPsQiIxUhbjKrV2bOVW4kMSxaT5pKYWY3RSk2nBP3Q3px8Q8Qh0+AAcYL499kTjr5OPw3
SZ4brzNx4HiR8fVi3q36iL9FlM5NNjBVZ68J6YMgUPBlLx8hm8UsCr/dYNlT3BDdDzGyZgKfDJrC
iCsj6hM6FeEpi7VuWbYqCfI2bspHoLgCNKfeIWKA4aXi3R/cX52fmh+1VRvFYhktMjGXCEOFSsAk
ceEAGK0nibWsq71eTtdtEVBxF+hut16ukIgb2XjDsPttqItP/k2AyhQnoFHiy6uVmhwxFO0aWnJ8
p7IngJGDqaMmDgXBY+Q95U4a/8s1m3xWdTkniWlfPTJfSDa9ekaRmjJ59XR5TwtadKqmV93cvReC
ry+iV6J+ov4mwlEkVM9lkYSqVrgZqbLTC/lpiQcUaHArNyu10LF23zOfxGWNNtMYs/tbj7+jKvhh
+whdnOUvby3CwzjllouLNyy1Jjc7C4/9jZP7zHsHKkpVKgsGXSY9rnKvZp1ea0Py20vPuCfsftUk
rkLI3AnmCqfqTXp0JxgsVPd8RnnYvopZvYKrvKLE8//e/cWsfkEGRC9znaWoxYIkKTlvHiT+TsAU
dUXek+LG+fYzaJDJeDdD+86fU2suMt0SqrKfrTa/d1OhEsWtGdUO0JJrZKrAz177yBNtBfLmImBd
s5XuY6kGI9u/RohTSUic/d6BdlTgpYixecMtovZ77YmAc7H9ZcWPTMsQpFLBPuXKzUV2tKce/loY
pHJhcvfddOLHXEa5cG2kooMN+/n9SzAZ2XAKZUw/FPi3Zws8iRbppRnZfzQUYq78n85RPrYPc9NC
bpsVC2a4cQuOcAPBnQEy4A0NgYITM1Jsh7hlN+b+ePA/7BVlirZcewKcGieTM0l79gc0zG+9NSQM
17thRe9j0aAFpxNVUAXb4EP0awblQHRWK02D5Y1fT9kO4DqC49FUmdDEUTtO+++eVfFgq/LIAhCy
cqlTHD8AD+R/GiSx5xZ3ykTzUXJY3BlMzB+Mvmo4m+hmg30NQE1/jspSUebxu5ynH9kd7n/gJi6X
d/w0qdurjbVQLXwmMbyFwwlY3iVhktOhuP0XyHJt3Rys1tevG7FxjVWDENRK8wr0d69/5vS5TccB
7z7LF4/tKdSJw+/I42ykNr8tdFQ0Oz+1qc12/7gQYUytrWlXe+nvYjUi0pYTEOvoo2qzqlQFDD5e
aV/++0hWzx4oeUpvQhPVl4y5K26zmObiInYQ/LE7msKVer4hNbQPytvEbVZGoVioWF0IolDDywv+
r1t8upJJiL3735vcaRI96fMSfkFUfSKRpdgxFzmghICLWDnZ+dNlAtvMq/ym7mEIUdIsEPiR9P1J
RxLkx2IvcJgkISC7bwAswIQQ0sabOwgO4B54kadleBZiDG1Lg9THOoYWy7mspNZuzPxwXS+jDESB
8OU14hUDY25L6gD3HhnuKoSVpAuZBqtXcIB8ayreEn3XIxe+aMj2Cm9inK3aCMEPrSXm6GxaEbqH
eUnqLkYsuuuy7kx5hqACrXZ4JbpjT9A/JuvcYsG9klqLJK+VIzGtwmVv4iraGdyp8arOSKF9VHBm
bBsQv2lIgX0PljzuD2WwU7qdaPIT+CTvIBmEWPjxhxoy7Q/xDYZfRycL3Ew1w7eCnjIAUSAKMnGx
XKpQEfuCtzmpZFFQo0v5tmMb9Tq22m+ZsyqheEL8EvXjo0Plk0QH4w5KqiyYJfXC9y3hJ6/4uR7k
UOnQbxf7tVB5Ad+uT8+cMQPwNvIPOk8xWLgGlJJFcxre3HrgT7/5nqZz/xY3dxYBfgHL+OkNEnSg
FQNbOjNyGURSs2A6+bkJvwndTJacsjw/x7mOfCyU/11F99B0uPRO5qf6R5Z70UT/QFkGY//fCTLV
EoZt2QTA+DSoDpGJULy6VevLaCS9rSgzAzwLvcvvTweSQTVxGmvXbHw0/w2zeMlpbclU41hrZTTh
ZPToN+z4tf93PORhhg+xedY23u9gH1Iu+Yv58pJ4t10pkfsV+uZc6nVHa6x/OB4vEFcFjjyCs3As
+qkTJod2lGNqYHbFnupNYZle9yxoGnqZ6+I3XBWUz7wK5RTqm1WYv997LISb0tNegtp5vy4IfQ9h
2Lkc6r6iiEMkfxI4SDVDUTvPIAbj0pbGse5RthVa3jOcGAJMK4i1j0cOZyJ82ylPqIzn+g8ClxMs
SxnOidZyTETIdbfhzEe5u0uvtoqOWTt5bEnFussqD7ABD5qnenh3VPM89xkvbb3Zhdzw21RLrN2G
BHrlT3GZkUWrUNSg1I69YKauBw71FvrlAHI3MLmMHqf7n65bKjQnAh0mHOikLYwzwnU6SQBTElsu
TjPOc2KKb/G7afsW1isTAeq6kkzhqtM1gtil0qb6YhuqjwL/B7I7PagAq1FVrXiJ+CFBPMtSmInj
KYX+2VV5Kxq1DzYKADtERpw8+f/9sBhif7uczd9vsHVcL0MtXTr8ESsdEWEGtRgcEv5tc5WutT8a
n9nvyqKT1sU8NB0kpDEASYhTd+kH3WsieZeoGA62BPxvSUzYyw/bYGlqIRd+9O3YECFxfC+ssSCo
k+OpBtK3OG4e0t7FeQ76mcwISxTUlOPJjXiqXfgYm3/XWWXxURK9Jt9CBgDpY3ocYWoAGz7icYET
u82gHXeS00NCdCZzWRsROMEVDcKy7/Rzl14dK7MCDeYDS5zU2WIS7fZ5RZcgl9TeiHp4+7W2a8tO
32Ry5Ct+wxByj+hIQyyViR2LFb6NksRNOnUbgrOXSjBPnA++hIEttCbWomwWkTGHCzb2EUaPawq2
GZ76mmjGAxviDWv9bfE5nyviiJhuCtTvsAPBzvfReL/pRjoAmYl43MlyygyxrFDPw1aXhA12OXHw
R9bfDO7xPYsj5HRDC5BI4URprYsLc80R3ZGOQFUym3+OUsuor8zza1qnGq89GE3nS32SPYvSXglB
FzQzBZUvn5R4ST8pHJ0Zt6DONlqNzjoehp4ON5NQn57it6WmnJXNtsOaNVSyK/maparLvazawmtF
8ERxH5H4rh9FmZy8ZN6EwHWhB5cgMCM8S2Uk1GOsj707Hc/ThvSybfZVc76+A6Oek6TuwpoMEdfW
Sq5FW9usdAEDSTmzL4p9ABH6w2A7+r68BR/28rQzAPQyb8glR2QPZvbitO1Loe1bmt6F0xxZhnlO
heBbueFSn8z2wxS+IoGirzcaRiKr8T8ogV5A/fwDpV/30BOmijx370uMsycaN8kUvI8PIr/yp1go
iLgPZ8kABhpdmxsqmfV5y9tyFJ7JtjmG9Yj2AaUbPgmdfdRldKG/ot7NmpY3qS1sHtWKZdQfjpmN
ZQXA+LmcOw2Hoo3PlLZSy33DCHwOPcZOf2xXqjdCVMc2VDA1BAEqPNJK5RQJo35WJdRBrgMTgOJX
y+KpIy756hGSoHVojtR+LKqxcgUoe+lMvohINPNRFNtvmHMqo5AG5Lo9hGQNwCetWochwgF4nySF
ZDmGFZl/Au1Jtu4oopP1DsFauC6uNUut636ODPXRoP/Y+nSDiHBWO8w/e29UvHmqLUBAGAn8YGAx
NNmVkxvX+nu2g2t47h//NlkB+Y1dFDKFcqw6eHBqXFLypUxGFkkutA80s9KqE9SyWy9tiIeSh2Ub
J4L0k0wlGsBPL8RIFYU3x8KJ0NmBpntTCrgSjYYVt5qBp1UDbZsnWbjHpS8f7PF1o62C+WhDtcAt
fjnrjABI7+LuKpuAamVYuFwltJHZS8BD5qyebvQDvU7q1mw8++M7QbnMX+AozK+t4iWzOpvZygLg
v+fcgkuKJEZ7uXPoCKDRKs+GLVMUtuIFdWyHHzOxE9mOPCqKUIYYo8KUwS/LFunMw2XV9oC3XaYp
KoQrmOPGBXbbib+w8CSEbtFtw2SvW2jTZgBNhCeke/4ghN/2u8bEl+5NuXzM62a3loplyimP+do0
VQBKUOVfWaIkKUb0PPSizhWWh0z4lhvDU/hl2o0dyj+0bJoqgDyOsOQ6KeD2EzAcS/sjQMwBZ+ez
oOi2zb84jcK5zlmyJNEHRKlo5NGLfAI0rp1D5jnFRVPm/oz0NGmrgTiNivEW3Zy3qhLONNF99SSZ
T+u7uHfGnH6C2qJBp9IC5GohVf6sze3Oa2rrCNbCGU0ng4oL0jU+6lOQLnmpqDkXFFq6a9wI7dCx
pNO7/U8F+J2d4aEleril+nMdq+jYX9XkMFM4wQHwg36OSnFxZE7jYDiYGJ3JN9DiPWku3Ec/nDk2
2uGKUiiVYsfQ7G4UK/6/VPWiyBkjZTZOiaL3fvVjEKeaUT+liq+FnymJpReTjhd4ly77NOrCcnX8
udvYKFqhsFeAEk0plA/WJUKR/FMiSEM3uBG2eY3M47YVKpjvYOEQCKmbhyGyU3r/RQx7eiFjGG7r
cqPFe6N4RgsSRjqNpT5BczICcnebH7i9UHmoCrLfRo73rhLPO22dlpB4oyrO9BrDbqWPGwCDYL52
zF5KpovZTTZnHSxumHb2go4G4NCqR7Y++ilfQEG7QSUnELtdDCXeB5c+mAWdSeYArODfQRenM+5N
+K+anPwuB5bl4yY5Wg6hNA5RpHJW9YQ0xPhJFNv8K1OXkOeMWECV4NCdbRiNu9ggJYo+VlUdHWjt
U0KePiNb4Dk6RVqnQoiYDGCt/AQo/y/EyM+6EfSBkuSXQqxcNuymlu5/7a/rTTQHiG3JYLlqRgRQ
giRqd3Ju3hJ1DgCl2Ygaklt8HyPu+nWdP7HoZIkyqxTysFzVufs+PeDYyzmZD467GltELAmTjsCm
CDQe8ByA8JSjumppgA07HnTIwEuSg7rxhI+s33NBnT69WOrE7h/fGaKzPlKLTmIfMyWdEEki8KxQ
QWRBi5On9J+y+bjJaEUbyCFu7XAAlAfE7X/S8csFo0ar5ccFrrr7pEYraNyvwMUEizfLhXfJVKED
37K+zgSGtEhMIJtMGoHbzMYHH7MCt1075ZCljMg1ww8NE6qlPunRJe+TynUTxOW1UV/WgnRGVmfl
JRom9BlhVh+55qFqwbgi2I/FE73Sjohtx2cV2+2RYF1e0Oi3iRGco3svmpJQBlngBmCPqB99DhHY
Nf7uzgE1RVJy0rrXfP9g5gqqDVRaCUFOPjiKejmBkYFVA8lGSNzucNeNBdW7L7VilPugVOgRT64Z
21DHde+qCtI7Tgro7rXPiGjEWmxRl1hd6pySr3zE0ALgYyUElFFYIptunoTmDsfAD9nOEInn3IOz
I6lveEmj3lMgVYMiCwFmanzBK4Q8/Gy5jZL1xoXwxXEcO21oxVlIjAgbpNa4oV2THHAd610kdKMu
RBjTi2U8D/bUcWi8DP21YZrvASos0AUEGuKBPJfpmv/LNvl5X2FevGDxSSsch60AF0Rckj17dTln
akxbTpvTKjh63BlzZJhEN9byMcQtC6XDhXNoWZ79Z7MHig7wBKqWpyd0EHoET+Tn53LceQ1C7zCM
1qtg/reCCPlPGXMbANIBPLBYYrvLBYyW6S96iw9x7U2lLW9+BbJMwBYofnHjdxNV4g0nLc5AgkOZ
7m1WCbExymJSYizYA7qSAPlBsJj9bEnfGkdVIb79SEX1Y8aDnexvmpEDbsVNDucvyZja6hlfeRPJ
ptkB1RgPZFtj4/HgZceXJC6SFtXk6RnKrCJ3+CQSPmaM5Lcxge0FKbha5TuTtb+g9Kf13TZ/k1sm
75IZOl8AXZmKAat36bsshRFur9PnCVfyrZ187aZP16K/QOQZYX5ThK6EmAlorjCH9YWDZvwecbfl
MnXvzxZQAWWwMbVCCvvl5M7LEbM0PRjLKWfESnpda4JjgMVpjYpEqDLzoCIy9su9D807HGltxIzy
QErJeSTsNuoe1eCRzEf+8RN08JvjhDedzZVOOJW8kpKhF/sopeFnibOoCgMQZtQ/+hp9Kp2A0EyJ
cZpKulyLfUX/ckGaWMhxunmk0D5w1vlESishL2s9CN+A+MLojuanR4IB85XRr/F3pJ1luD+KWGf1
Ia4v/YjHlWzA9Wz9Lh2jq5XRdc/UWrfzE0MNNvDgXnoGhcZaTaRX9O5e1cyoaTCFOHJ+DzmKXTpS
w0rUwewI50qRSH+IU0CMOswG/678RlqqbKlDtpZ8rWC9fdKaoZwBY4jdcGJ8SkxuGwWisjYPaMsS
yFgCnRiPm59QoI+L0WAd+IgmCr3SgCLa9QfoQ0GXAJPKkqkYqSW/BsWflKt7ZI2iRZa3NyCng53T
Tlw0d5uqp2YyEBjStqqVo09ub3VBMeH78DzoGRsapPXZkXqjDsyj64FSsdGqGZ9sGjYpmUGdSHzY
szPDLa1TExUc0RRzzlamf14uAjvYcvlj0DIQjzGEqWJHgeNSePZE47lnAdwSKA7NLarXHnrurK4v
A7QhCIVAKAbWHceOPZ1/amv4LIp57H921Wpr6gH0zZudlw7o9A46+aeq/5UdQhIKfAjQ6yy2nogx
hPjYVWtZpMYT84Q+ckpgbq82WPuq/f1pLx4m06kwn/hW6KYk6W8gjQ51OnYkb+WRxqf4grTcAb9d
nHXmPacvnF2vzviftJAKorAnY5q81m7H1qDWPN7vBK9PxFR86OP2wb1lJn+7pX+XHzbMQ5CxWG2T
ugpJC7k+amw3l3VoU532jelt7+UDp2n20AJyD/RRhyuzh5JZc/Wmy2b4k2c1jyFkQRuoVmGJc32E
iqdbVvivRzVpcejSUyRX2SODPe7SkaRCWSllmpvZvH3ghMGS0RV7nFed2a7R9k1uxIQtG/v+/QBj
9ttZp0lbcMcmUP0uRFmXwwRhMACvsfuy1kXtRNf51bK/DjK1ND9f3m6xSvSvywfrtoyH14P0ML2q
pA5OnKS3zvNEykN2LEuvjwyAY5dlzXE8PVCibYujXysKa7Zv/fwKjDOm86JUpJiVNCrtI/KU9FiF
bfnZJlrYk1Jm7KMmW/2oN+hHZ95rNzowgi4ufe/4NSIunNsCEQtBPoe5S5S6OouKqqTJ5I4OYfzI
lot+lQyKUFS+Ds3dSnRk/ex6WlRj5kh+jMBH43+WBgxF8Dn7540oGMI/nGT3aRTX4g8duabagYb1
ZwnBr8K9RpYGURetNtGab7UbiKZIeV84XddjdQXipSo2BEYgYMDgrBifGhCW6gLcVZiaPWKfOuwE
2phQnIHFKTgmzeh7YxHF1mkrmdLnbxPWEPDQz3XmKZpxfzKO4RkLAugL+f3IH1pI4jMyyWFEPYyy
wSrkbUzfU0CkOTMiu39UQi28dslblfqsYq2svHqDZJ9PYt55NFBtr/5cPnpyNGF/mKnipWitLPtM
gAARnM4xVGUe9x4AOqDe1ojahLXFnmcbHMFzM36fZh2Rygg+W0wKozGnxPT68Nsa1jYJibasdjXZ
6UMfJciwoLdfoKSSa4xsQOygVQisTpARiYEnHbCFnEf9+1F6DrRWkRloqh5YKX3+N6H5u5n7Cdq/
omaNccwZn5Y1eHjHgIH0U5YWYoirDNdmwc2rT5mGuHw8M0TcjO4jcwC+cA67QMtfS/f0Ks4vVIO9
CC6SW0f6m6AzwGcNsR3W4vXd/NNqOWKUu3kJysk6fms8G3UtuTmxoDpkGC/ryF5jpnkFzGbuAi0K
RMBydfZo2JmDXPKcQ13y3YmhXHy6ousFHREurtNfZqUt4Wl/rya2DlfbgDsWyZ6c++PF/t/+Efhm
j1EdPTm7sde3Y1qzv7kcBYUfuPLK1lRByjQOXOx9S4mlDBOXunC++XcLADk5Aru9zzOXbdw3BALd
5BZjA6GAkxL1E7Bnv/iwFHoD8NotXcEkdi4jBLOW8lXumCzNvKvFx+izaAfagEWMZzXv2I47MfXf
zp46iaTt39jjmAREEhsl5uAEsRJc6qnqo6q1fH7Cal7yWIjfmZhQRLZI1gUi/7foei8WFgt4BLm7
7rOIZHeOspXaXYXlN+A6Dig/GeOX1/WoW+chLEuIPQOhgX8y/j0ELxgppU2u55CdDDmwfhYsJZCk
H9Z7Jx/FS8OAY95WAwI59ssHE6qlDGS2bQ4zYyVjH5+mGKnBKDr1vjJOJF8haV/cwgnMOD5y11HB
eJvKwfpAKa3rxm92w+i3mePRtrk2zqQdh46gc8x0J2KR9T3fyHovqQ79HVl+wb4jEirwy/KRUd1Z
15rJxKnWFrsun1gGnh8OHVDv9926xxJHgrUPJxx4JTERLpcW8tKtF1/tdlFHG5bIv/9gOOmr0OWE
jF7NWH+Vr7+tNxXJKrS/crr0MLZiKRV6cZnUhd1O4j3mmqZBbjjtUaiLjJ9x+cisLxdbeGvJZ5QE
ajdGcvrtn7sGjvtNibDz16sLUHmLrEggE4SeijxaYEr5YP8fgtagesNcGg5Ukqj7aAuYewSKPPq8
Z+JfJQ6uP6fpypZhGv+JDlgQx4ROIQ/tppcUnTo/Sv9I4BjpCyPhSEMy4aEzFd5hgNgr/va3RCDK
7YQeqSfJlAdGtqftWnCOhdwa7S+drF6TacnIPn4xLr2xYDX11qWpbS7bO/MOJvb4Umspjf7l0gmP
MMW9VV7nPpq+KqJAA6NMu5TGvZFLAHahgWdWymcw4KKqi4+RzZ0SYTIfSmhYBE5dsc5WtAP9TwvF
Si/A7UzA46pzOzg+7YYo7jVmhSiu4IPl6vCe8NNW80M4ePAZhDZkY/yeWxdKH40MCMcvsgEI0ho2
AcnYUyoUCU3FYnNx8kyJJsf7qmyGkgmuBk1tIo4yODO7cAhQFroWSMHfju4wxdESNyUjEH5ezSzk
QP8HoXZCHRWWb8UffxSfZ8JuDfvk8dd7/IlKsakBHRTT+3F81rzAYEcewSOBNKrp3qzYW+TkJgKt
az/+lM5q5tjBjIpObCBua++G4I7Xbf2U0vFzLpOLvwJ2i/yp0mQ8fqZGzagjAx2AvnIz5ygPaCy3
nE91QU0NuSLZ9jYEndX72PEcw7pJJuhfM2NgSYMRMlfA1146l+l86lPNqEc0jKkvpHYMWHhR0SWC
+oywnAZWa6znizJEwWx3wiCF9LVrLyeEM5nEkASgRknx2INXpsLopvv8h58z3MYGGtQO7C3nEGwi
0+PTcS9+SahtAmGxDmS5K4An77ohr6KBrcPLY0CriYCJUzX4+Q2smTOX74fWmZMA9uhgmCdaFCcu
GJSm1ChZWxuZR+cJ+/Y6asf0c3CoTy0HXJuP2xzPcfhpRaCE3uYkM8Pt4Xxdzh0Qe8lFJ8oeRSZw
2Tc5FFB4tyG70r974SYUPT2Zs/3GpjC4RUt8eOL3gDaY0kjQ+8PI7BaRgik3bdHDcc+ypCN/rEsR
fGSXhfySpkMDh8yI1sHnzN1/wc3CAJjLqfs20aibTXn4uf2lRpClf+rg/z5gOA8lIee5zsQzZj1H
XcyoYXXN73y2W7tMZ58jmpADa4woaQ0LYJUCZuJq5n5XFlTYn3zxmWJxAaNTSvGJUsOFFw3mGylM
pzXtuqzkDEgaW2VmAI6ksQCqxfHqqyoubHgBImMdl5KJN8I9LWA91uaTWR0m3hTtuAQD7LKPdbW7
Z4XLMqWuGGysyvxuvscXyz/UPvDJREcsBQssMM61zkEts/5HVKl/2ZK6dg34zUlSkFjNduwgZ6ih
IxPKu2Am2iVf5O/gFrPrr5qwRwiyRmChq2UoYB+CmneZIvGJra5dX9E4rGt+uuiQo+RHk4rlun8O
oZj0SLVH9QIA63fWQpiJ9Oj9Y5mIpB14IFAF13yYMRUv0fKVvUEfIIbyld1OlfaFJ3AO0kiqyoPU
8qg+81mkBf27E0M0BV/MngO3XpJy2ikH6TqiUKz9Gw4RSo8zkm/N/BVMrdWk3LDNnEbgoqAkDX9h
RsHGzFsBEdzLT9FdSknvylQUkv3RbOSY/HQiiQbVZJPdt/r4kTzwyM53znzsFA51ZFRAzwAsZjwV
i36pKu8SnipFvCkNYSYkPLYSqpsxY1HKO0U1cyTeQ7/15j/U4frNq+FJ2s/f4jKEahgSPgIwHyQk
yxAnmm4BJkiN5d5UnCwX8veXbceyFFaJIKf5WP16PYjtmKiqN7BdzihpIckAsHzxiB/Sot3hNtsZ
GoD8GpFgfcoV2SbO8cy5mVvhUZoDAcv4P0KLyDjgJSG62P/YQbPcVnuS8u9lxmGAHZ/n8b4JK7dk
+8ckz+l1pU50hYcJ/QHCySqf7wRHiHbw1qLGqkeksG1NDXiqhC9nsgghDqXR2T2WrhrLiAvbnJk2
wAFazoW1emUfZg2eThgi7/AVIefFf7/195Ay/DE1PlnXjmgvHQ5V9n8KMvAvOv/b/dJk8zbkVTO8
0CVveo8+ZMIFc4fJrAm7emF2D8HIJ7IbpqLTnz2xIFuLgeTr/+V2W9+UZCKtABzcIAC3uSNoRjJt
WQnbCJoltRoVN08gR2UfZnrkNd7diDjgb4DZ3tPaSuC2cW6aC7JPLNx5LYx3+uBTP9OAUm2AilHw
64ITA86NIZHbPEOKNsp9NdXXaq//WC6i8kgPaMbtNLjqD/1In1cdERBYh6WLcfWK99Vrbp0xJwtY
YbekPXnqLoxDdz5gIC91HgeT92h8jLf0l86/R99FUvUuj4BS6K9InNxvGDxhOSB5ubc1zfpRPU5n
pylbcHC475kOiqkk7/ICu9UvCFliGNKJb4MiPwOXnZc6mSLpezmWO2EcLu3aftzuUmSOWKGBIP/W
LIoA2lryqSA/x6gshCVBTAHYNu6DaTLKWHMHQ4jKIUQksz7bz0DHoxMr0K/uXH9ka6Pnodyj9u9A
7oTCWbn1baxMqCCJxFwujzIoQ5oANlQ2JxYkemOg5SZbXO6JG0sPGlJuEmtIqHetg7Sz3hOWOjyl
V4SWhbwZslqSg7uQJplQnhufJfvgQ6amQSpUoDUB+/h8wL8jWQCAC5w2rEaWLAbSi/RGh9HLLRD0
7eRb/dySLYvpwYSDwJG6jm8Pw1VLZD/17Y4qZcXN+Ha2tufX2gGXbUPHCnEOOOCLxVVZSWoTULDF
prl6bK7oBVH6tu5IvtTJ6K5zrCvsJeqCvOC2GQDe0X4c1dFVa5/JF9aXwqpORY73kYTgxfJ78sYx
+iRx9msssKqoMedspFnJ0alUWUlAXtdKwyEIrKEaXydwKnTY2gX8TEh8SGb76ocZXOyCsElH1uqa
r7g02W3BNL5UTl7csttWfK3+T/pCP4hRSH4A72TXQ9lv2Nxu8JBLiQCxc91+13IBAnFvJnbIUyWR
AzZvuuxFvmw+Ev97Jo76K6jKBnLJFWkUCJ7RwgsYM2YKelOghw9NvZNv46DJES2CukTukMi/jupw
qg9K8X/mo1750c9i/W69Q9e4gJISsFnJJWkpKJ9WaGXQyRpg4476R2GTYmbSiTDI8lgrtBTZTnyl
+LYnSB/P05OCSqG+Yz7UAtNo+mvMRZfBB64RWoqAj/yO+BLhXrY1nSs27XFLAY5ENbby1gWPp7S9
hYSaJReW7pLjWk5Fp29PvCwQpFQsZqsnUImkszJv3qrTkQMQdTAhX7liXknvNyFUtWq1FQK+MwZV
SxgwyAbpcc4yJTkyOm2yOUaSxmO9ON4e70JppsYzRzcrIR3ypp50OCL1RBbq/ysi9ZGwsL0DKx20
rd5OXTBvmihCMShHcFpx96W+kbVvuYhhVl9jQzHGawMvoxD5wANRVrRd9xd0LHnxoj8O3kjOHL0D
b/paGx3om3zcEw6n/I3X52UetEDarGqF+B+tDP7un0qdosM04X89VcEccf+3+xItbdRWtGpjkokz
IsH+B2D3fctE/LrjsNqXJbFA1364yolWGjOtLhFJE4u3TBjdjT9WlA31ZfD8owj1JjmuxPJUxW7E
geT6HdW13WFSVbVGHoqqpxGXYkFPUdOrQu6WyYrNs+9QUHKSitIjKaUGla1NmQGe+Fo3m5J2upkC
liHRgsMhwNTPAaM1mNqxmy5QCD2POOnMnKw6S1eVMQmFlTzHJsrPzthA7v0E0H84SA8O7ueqXzdq
vXK4h4KkKm2pRpe9cVXA+RL+fah3FN22JVR6pdIWqB+M/i/5y+vcMhqzW3neWi+oNRMRb+wiXL7Y
fcZYZsqdIup2MjTg3MS2o4XUz4r5PoOhg41nngoiGPfhwltqlcKkquPQk4njjVG6Ph4mMsy7Zlkc
NGy2HrE03iDbzH1MHC6tcvtVEShJ4Gi50x/7I09vrl8O0w4ifqOggVOeBRT6o1o6A9juOOxi3tg3
dzCJuK/zw1togW/JlAYXZ2cyky/rlStsmYJMJWtbtnbq8fVpUi4Wmv5w1K7swhKL/42H15ej8tQj
FLQCGoWUc2g+OqhetQlgTMP+cSztwd9iRgDjgxlQt5MBs2tRWev/OucrD6kj9Wl+V78pnjOx6Ylp
uNfxvtXRFebNFCrYGutEheipdWxm3qWsbvxAOw8TNGExQvitku0HR1Yv0Q732bpEYH5fLqA5PXMh
Hn/NwQZPfGFo2xGtD2/ifBb0NLKGYUKhEEYxFtl1QECB4i9Vwuk9nx9ewizx3tL9PlgvMz2HEPJy
3GVr0Zcmz0YLGya4W9fOzMOSsn9030r8Y+igBQIOG3vl12cxQbIZ0lH/HFlG6RTS+zGCtynCN0xQ
wOW+q6BEaNhGhSF2GJPPJ/OdigWpKBGdPRLbRY6a5SySgiQM9LWH8Y3VjBiPPhPTTYDvN/4G8zhe
bRC8RAJnJeRZcpUc6iKD8QFOnAMOpfo5ogfCU/TXOBXfxFgxzQGYx1G1esTUlYU+ZG2JJLj8ZtBf
MKkjPVhVjIHs9qSLngoMI9MAR/86DFNI30d4Q3WXs0wT39oBajGUEjylENPkdM9HN0Q3KXZ/zqQU
+ZEpCHFaCBGrzsOpHRQwAE4c3FiEocxDSAYD6yrJ6pE8YLWS7vPfjyZp7sdveIZifI9F5IBLsX5D
4l3mj0SjSFqJUFtTCnD/hkJPj9rZfkjkMiM/uR1iNxSh3M7PnQXXsuw4R9B5sotLXq8ayWBsXsf8
DcaRRWh4EB9/6jMe6nI4gCNjjC278euBLbK2FgDiKVr2RTQ89rpNthp+/SPv2VdnmZ5QGU932IHV
co2ZvpwJ0NFV1EMFPBc1czrWKRFljXo2wkaBeera52Q7nfoE50Sr24urktdKsxm/LTm54AkH+FoB
L9wIUeDv3FknZV14mjy0vbLF79unYnXoIqrSMCwQsQYxxLyUiywwc12gShiYtjtXeJZKBV2+y6za
hBXIdQEaG5svkr5tEJUxMHx6wOvYJDso29JKnnjzMfHfvobYoWB8gCOneSs8mArS3bNCwV8slJdE
KthMv86GVy/m/DyEUXX8xYo4Yd/X/kTCXKK5O4dts+5rQfKyDfuYaG/gMhRGmkqrvpB3TzqhZebu
hw+hkh7GqCSJk+rw5wVTvHG/9u9aYMyPn1LmWGUOgRj2P+Jc0sbz0P2LOGa/bqjX8WjLBb+jePqm
pyLZJX9Y+VcZuxDAw+W4geBa5G/FFIGWb743SaYn1eSpLtgsvSmFESdZF+ecUB66LDMVGBl87lQi
guKT52H41wJavVZv+fZjtDPJnwujcqe7rdCF2ZsxNve/lny8Pb7By+1h+20P7Kb/EUmXhYhJR2Lu
AFaqaJZfXVZsch6BJPVZQ2uq7rpGLWekGVMH4DvLgPIbohyhFS6DJF7iPe7GcbacieRK2rKfqVqy
eeF4s7j2TKcI1QLksH3cq7RzJg5ISRlM5QvHE/3Ost2dbYbelffA+0NK8QBwsn1RnvYpVdQBCWKW
UfX1Mfh2wARouaT5y8o35cJiAomSaIfgnrIN+DQtiESloXBxVa8kiF0EwnwlSdJ02q/OpnNLwoAm
0Qpi3V8eGvqToBoXamPZv3oSFfjVqh00unpaSxZ5oPfqA1vyA1R00jwx5X9B5AbxNrXdG8yQJYbV
SpYw71ErcMGlwOAtiB3+GCFedUjFYukwpWiQ7VGPbHRg3Are5nvmTb401J8zKj5bP5e8unL8wZAS
oCLdVnKrh30mDQPYD9g7Y0fKpUuZlHxOWxQZMSD2iR8zvtKwilSo6yNYJCNvrxVt6a/TjZH/7JhR
4lkjjav0Kk5m4tAqiomKM0cvjT6Ah9QIN5OTfWQITK7e5/ucVn/o3cCxiNRegoaXMNUE6I0NvsSJ
ZC0klYrbF2P1Jsn61oV65x+gMizpvpLGCxKnDXBMJY2mRfres/RK4qmHmlOZVJebei1jBwsaZRpq
VmhtQD89iKJLRY+nBarphGAY/rJdpEd5RI+5ruU70M39yztS/JitmW/lnfTMizbAAUTbp07e/loh
uL80fffFeE2er1Uim8uk46vyTMEj5x/eOqsF0bDnKNFQ8epxrL2V/HWK5K+Ffc5loVxneXVABI7W
gs9csqbps6Akdef3xCTfrrEkhyjvRquk9syAJpJBy3q1HEStcguaKkuLzHzdOwtEQk1Wbe/aWGG/
Gyj+2wh+FLZrcfQDN0yVKDL/67+E+VMgVUay8EsTGoApdN0jhAZXm6jsk5+NTq3/uIQ2KqZzsNtK
7EES6TNDGM9uinAy0XXG+Quk7VpujBy8rUH6BnWOEB0wh446r0sp/Bf15nkC0tJa0SYGdkkHYFdn
SsJH/MLnlf/rlAfO9ubkil9Y4W201+3PQ79HLxXPJcKaeHZGLqv/8tt7LvsBhjgNS6+0XfRQXzbB
Anq1d/XML9GJf8lK0b7SATUWjQGegacyuqMJv65U/DN3WJx4mNg64cgm40vGxsETVeFUWD4cKN2C
m76pE7ztxQyJBJqPitzDXCk1wnr7j0+yNzi2NPiWK55QGubyrtenesAdFqXvywHgjptmcR2OHy1W
cuGa5WkCEQ6FTvLxb2ia3o+LoCuiHHg6utBEnJrzZMmPEu0i28400yygmRwPMeTwc8aA43DemwSL
8Vdkmoodw52RuPkczricZm1lENylfYBoy8dwIhzgTq4cct8CNlMaCth45z8kKSbDSnG6NFXTNf2A
+Nv8fvxEosc1QroRoSUr3RQ11lyKq3DjbuNgm3ohISVYD+y9LkOt6COqyGL9zrcvqmTEAX+C0wz0
FvK6UpwL1zdfVBqOl9e4GWkbyIdFLur2OblYZY3wZKd57CeET56Qag9P2DDajyFHsYCDXF92klNr
vNxluAEfvt+KbFBc6qVsZYWeeH/TZUHBq1A/6sQplD4t9iNNqURVA9xcTcdrkxpTARZXMEAUGPqY
U7tE5dkuNHAjgloEIB1zH/Lvowbg4hbhXpTTxBbidcExcLJlJR5zH+WYMxvE+T07XB4ebE0q3iGm
Ty9J8XofN0NT3dZBChdIIHcTIirzwYPTxyAh9L42ngC59GaGVE54iYTd+jtaCLD+pNBCuzvEPY3V
MqZo7QH4FVmRRHqudvPrdFnTTZeP5BOgSoxhHm2Ic0+NCk3kVe4TofeF5tyFdqiQDyXKoPFsNUps
cSaT+B9HSQvJeljW+Nw5QPTDxufPSNPwoLA9zyE1zZDRsz8GL+mWyqWPQAAkVNhpST1o1fdrYgLh
T3t+7hFarXNJdMWk+8Z+1FM05xKDItoJ4JG0PoC7XMBm0QF6GAA+H9H1C2uizedusy6nL99GZvjj
zyOyLDNf5fbNXDtuXtxpAdetFg88dvCNguH4SNv+ubgluvUPG0vgqlkC3lZaKlr4PTRT9hsTFeqT
ttAITAEklYPfNOuLy3DYP+h6XacjaKyOCtmP3/nrhOH4E1lyZhSDEuMI2DnRYZi8hq8UlxLZodiT
vBC8x6RA+oNVsHMuxu1H7IAYX+zZwtc4mYeY6SbN/cONr/U9w67GsuoMP2hejTZuRGe8p2S7i6Ms
aChQnHqp3hlgx6CDrGFTfRSDarHWo3qw6dfpyKb3Q5YD0U3SxviQQjncsYwHJSdJIYs8MV3KtlWF
GIKc/xp6zAtgbkhNXHZU7jBlFIdjj32ClhqMM98acOaOVNNr8WjyJByteN67elQy9J70a5IXnZ79
nU7oOxpA+AsN3iC8RfH5LZhDOBClk272x+Io+Ho+w9zvUM2aHWBNc5nUbt9h85kqSRi0q8Dkb5Ck
UjFUadmeKeo9z1jKtvxZi/JydK4Zmp+ZeGtltcyz3x6tMISo0jNvrtXQEUMoS6p65lPcliLR3/Ba
ZPJcHOABOmiZACgk+UECXYMF0Ab6r34Gn8se0c0+4lcHSFfPptL839+GGXAzaGL3FV2ci/7LIKCo
S/b315WLpozS1HyxWoE51auv7FbFtEaOxWSDDLFY9VETt5QPOXvefHrPgs1n0d8PdK8Y47Xp+VRr
7gvdkdJkK4JrDLbMI02hUW3SGFrsTXaBG34fa/HFXbaD5Yj5U1GhyaeTN3MHRveD+fWw+7RGqSHH
IWU2P1ESF6sMh35VH6zQyEdGyFicAgw1Bq3YVPSGv2blTygZx4+hkRFi53pqUVlalknCMrhLcabp
a6vQK6WDveziRwHjjkr440goxPQkzco17uKnJzmSk3dZJLvfaOGF5DfFpCaRjtR6Nm6h1Jw3qNJ+
ZlcqRRRyyjE9noNJWAOp+RWlEO5hSWOMvtophaZ7MzJS0ey1F06pb5z1nSRBeLKxKOpJ/fzxlTec
X1upyUzhyjzjQFs221HnSxGREeLsmgp3C4m809e4li5RIsc5RIpVnuoUtQ83Jbel5KJMooO7Wfmk
CLV3UB5shxaj4QVF9ddnETZiMDyLiZjaa03iFjKl11elZKO1fAZSfeqji5n02zPYDIE3+dKO5RD8
mqrzklZPiG7Y2e+BgQdvBxf8MZ/RQaz0KwFHalWzZjV8Rm8S+JcDzHEogikCZkjdPvYeWEtjXNtF
JYPdu0GskyKV8iBD5OeVmzcVwRbp1ebzz7P1w/j6dDwQRhNIIsVzdIRcEpJqNfsTZSqgceR70wxz
TJ3UXpz+X7CveBC1jB2pNX8Sgu/DwhGtfPdaEBe19KkFI0CkfPWZgUym7Mi/lszYgs8udhwvZxN8
CBzWr0/vVKfAv34fJtQwtt1xcmj9E3KB4znNlcY2iisN1zERE6OZJGkfbHjDtoGjDUdS93JHWWWv
C9KVWw/tq6wmrg6Vx+E5X7PRCwbIyzjT7wT7Q4kF6xakpajsMdgru+c4MAFbyQxS3depLZxGf6Hs
pAXihE9gDz3r1qasRfyQkxTjG/NQxzaxXaNV+ZABkGXwuqEARurYHjcMOn2rVisA1AzqSGjdyjTA
46cMCwKu49DI8YUfsk04V87P4Rf1FB6PnSHxeaKV5i6RA22xFNB8DeAzHwB3oejJeG+KB6swXbgo
dcVjjTxNt0rfhYYVBLCCLj+Jf8U9H2Tr1sJT84oa9fsAo6CbQFwMOiHLSzxt+5cXuer04BiUFsPU
RbhbZR8f7Bz56itfh513jseVng8DJsZzpitBQcjJmGOXzSQeSV8xNvxjSzCWQFxwPlPqkSie2IJx
LBqhbWF+D2Fw1olyp4IAST5uIypaiBH4gNYmR4Pijui91AHJvH/XZO9KSE1STd03HVi6r2L2svo9
nxbnbZrxVsLSd/FRbwwUi8wGqXL1ODhUOJKyFi2bUa8dqGMKeo7TLM+MAOyFnNUOjDhkKSowX0P9
Mh6QlL4hbEDdx1wu6GHx8xfCPbA24TWfYf8Puyz/zRaCeiv924mo9LTn2y6FKlS6R+X1PnyyHaJ2
kA6GkVR6BP5Pk0gv+agC9BfH5WIZIyPG4o7CY2UgPG8hImoK68V3o9+kYW/KC3/7S4hmKMpERXae
L5CHeyt1te+YigxkEPWPYxCsshYhqEZhtL0pCio7r+YNwg6izKTSM+s7mGBYFa5kRi8pS9wlJduh
s7QVFHn2ZWkliu3GAnniLnKkot2yxAcfosy080CwUFr1T8hc0v673RjlEFvs5CZa47h+Drd0eeXb
huFSUolsgjfrkjAJL0zOwUiVfd9gm/wUH9Rzh0SMTKXY9jOZk/ZdjeSNQZMf5N9ndqVHP5txV6zq
AWoIEqFDGMFMvdTqeV7iXOvblxHXnNmIuxOmDJRqX46olSLlQDsYiz7TEr7sSI5b+hLn2o7Wit7G
GqAmoEHtP0IpxgwAyeQXhYX1Bd5wGHsbYRlziWzhwNqoGigwzMI/QR5XE38MtkR1v0wJ/o1k3b73
2g2MQt1WRmSs6SX5UABN5ogjphwlNedc+scD2jz9lyaOMihbSMOdQ7xdd03jRZY07hFmS4mSnub4
ttJ4rQzJx+zBQYGoIGKlZnmEgSM2C/ZuM7YTmFgCaOam/EKQoqb6hgZWoKhQFKvfbLZHgNA5xJTM
4oTIG+MJuSl1NV9dyPLl1JpWIkdhzj9e6MQW1M2QfK3AJLVgBAMdzIBE0bcHmXILJOf9yOnwfAS1
cmmq2fS1WL2i83NrVi2jdUgWS/qU8qjFfXK75iG8Kd4s2LATrXpzybR6d/vyUsgHQAHbQSsWVMTm
M4ufCqjNueW+k0+nP2ukZbnEusuIvqZTSKTABvC1IZaFzr/euFa0WCNQqiGffy1N7NQJjFXtLGEh
lIF/WGhPjM68HqT0rFSrzCZjMqnXLGZ80ZaOpTWxUWlNltpB4H618CgKQ6mz6MVGoxvZWYloantu
LyBLg7HDmcfoyDdeOScslN2SPVUwHhTgrUojykucehOaU6SeXaV4LJtlnO+0//zso68YaFNkFuyd
Qopc+eaDj7MC/U7ASQlPm4QBtNGgN00bFns04cfe+vRAdZ/9T/qMdqJFtFh31CcRVNXmdrDWKeq8
gkq/sxHytCcpu9Q42yIAxUne5lHyHZVj4Z7DQzOEA+5sxWomruCt0aZ9mxst/B1MXs2Zq38rA+Il
D1A3gWHfb9W/pcooFhP97k0s494J9D6/H4jT2Pa27IY30rdw+oIFf7v6IjMRARzn9XbVuoffTwPC
hEZqMdb0KFPBH5sccL8919AuJWN3yWHMRFZl2JfeuueSsXMj7Km7kuykWdzYTInkjhwiezZBa3GG
zQ7DPml9+hI6pl2rpwYpNKfcNaGllIAUcJNofDddnrCg/kbamQy09BJj8MZssNA2lXNnKZDT4tTR
PjVnzu5I75jlCBraE1Yr7H2qCTmmm/uCc7hCH4qwB7qlKLZtD1L7rtY2A8yssmYdEewWpXjq732/
q5yYmuOwiHcXuj6SKzFM2WJzAB1bxuMaURU2UG47nis+7dOfqN7TrpN/7XIt/64cK08gTgpzV6Dy
88+PyJMmnRKdmPGKQRH5wAhgpPHYux+8DC5mWjs9UBOqlnVqL6niHWUnnbqHGqAQ6GI9nuQwKeM7
FZPLiHAHgAOcMKLO0uDsbCDrnTWEFoy9zLcfAkgmD/dfwKW7c/fV6ljtIMRpKFPc7xo/qrDrOPD9
4UCc9mkxKWW0apIbmDcofeDrKSCqFNFEujWhCoBG0w7gWcYnHVmLcsv7ozco6IXW+s9X4fA6jOTX
MIV8Qh0x
`pragma protect end_protected
