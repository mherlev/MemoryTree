// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:52 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
AJ/a5sx2ccIv3PkUoI2cwvaPPbeSUxPaZfWaZcFmKZiNWQup+H+dsn0Du8p/q0Gg
4e6595KFroc9tiZdIju0kDTi+1a4HWNu2k4kzCT4hzYNHw1PfmgokmnaTjkiYYbP
ftd0KnSZEhAS7TvYFJFx9IJ1htZwW3XPgALskJ2CN5E=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9824)
GjH6RbWq6nfe2ECSTmZLrHk9bfHBs+uy5LMLcDYMrNzqcZaWO9/OclbaMHIuAM8+
ROqLr3FR2Ij7WvcVqxYaYZPpICI42xGKjNrrc03F0K869th5hDwF56IZPmqTn652
wQ/pNDz01z8PcjoFd6/JQYrNOuRu730yqdklC4277BKLiiTnbokMS8kEDhz6sljA
ETfZvvFQWu+oa6SiJJCmoRkcpZULxeMhUJTO3ehhA58fM+VKp5TkvqoS9h1Qjxar
hAbkjNjPRMgopm0CFigQpWDRAJNlOq6J2vo90BLdrpNsy7T8ZQlNbpr3fpfy6x0i
Hm/wTJ5lKi8T74El7mUipSu99D1ppx6qW9XKn/i5DfLaGhCqqqJ1pSAGKznQYw7G
4sA2GTzAj5eJfzfqKfw/ElxX2g9RvyO2+0w0H2nOG3JxxZWgI2Ad9u8UtAusmYmn
pz+EIJyergktE3GfWrjJzGfaBD0D2u/HOcRmGkp7X1qoSKZxVm+fdKxCZpOO2NOZ
nVU/M4XqTjDwC+48t6h5tRlthHF6Y8hGGD75Li+jVOVtfMNA4bvMG00ebERkBqfO
Y4mcTh7ozxHS04Plf2YbsX4IVcPwMwviQoJDNWdS1TYUUkRC+QnUgYoGqUMXA1gi
faxN+T/ABhvHBKLztIm/5cJmmIGYHyWr6YqSNOHPgdHUeKtSDRIf1o5iVPClsQ1N
sa109y9pKha4wCtV8vNCtEifkGeomDmQRVcomEcmDp5x6JDNaST0JN6oVzjWykZi
FC9wMXWO/pxngnG2y4oiRmbQrLMK036qMbOxQoBuTDyprK3VH8O0+DHgq+4IM/Os
lhENxHn1pFVVg4JcjYbibkwQ8oQoswjrE7g2XPui7LdfnF5hKa6mmMsfVu07fVk0
EZcheMil6VjNKvwWV1SkzWfgyVOCOWmHUwdiWwiM1VqfmcKjuJzJSzJKfsZfiQlj
lJqzknroiRbmT4/LObs3NULV1lygg0dUnk5mblDwYZtdD7jkXs5zHuK58BbKf8fA
pt9z0EiqUJtjp86zVRK0fG3GehobJvgbkVY9MBoKhyAypdMA3nuUt8f0ezCGJxKc
b2HrpEZK7P/NYec62wS34G5uPiNkg44evw2govn/XV6ic1yWmE2U4AN+y4zdo6w2
E83GyZNv5THwloWuzYZ6Nz6+yujNa+l9k8VV0ZyddF4rBCgQCl+rn7OkkuD1gn9T
7Qd9KR86auGPX3+dFgu7a7JGRVGYqEnGE7scfJQs2DYn8U540HB2YCFglnKTlcdN
lcrmbUdvFurjKFfc0/cp6Lr/HbsaqamPBAPudNQgrKuofGJ0gKreZ28qu/G3G0kB
T0XSAYcFz7F2fKMhSjsFGD1r8MYzkCvP+Tlj4xB6HqWHtjsJ5MUSUswwqePVVH+3
HxPnsWfg1o+EdBdL0XPIMB6pE8SOVKSXF9SlQIhJaeXY4fyih/vBMRwNAnEXJY5G
qiPu2XfkZDxgc66dyoN4HCwa9EDfEA9sLmOahle0vN4LxgIcq6t38kct331OVLuR
iTs/GbE2vonm+BjbPb03Pqcr3SbkPJoDEc9tBEf+RnRdMuh+7gdrf9ojS7kcPCqq
beGoBGzLDtFdAcTa6wra197yUP/WbWagZeWXoGuziyo2y5rJ5Luq0Mzzsdsl+Xo3
ApJDeBFy2E4ZNj17h9KaDyaqAniomvFg+g/fFcBg5M4b2W2HzYTFr3Cmuidmk1a0
TWXicOO8zF+axLFBJvEMP9oJMupbuIDFvMFgiCgjrZPHUP2U1tB6e8fcICTLOTrw
N3Z3/Nl9WIq44kIOwJyShF/6Rmx4TQQTYD0/IadbYJrmDT7BcGMueZnSXSuKtD1f
TSIKK3aUXZKcc/1Rg8WNc1r4j9QRUrR7iWkNGmi3hxagMRcNSS6EitKUfyfbil9c
IWSeakl2imIRvN715hcj0/YnFgA5xIfGt6nfwa5XpK1YZ+D7F7ObNKiadqa/M6EX
ONVg8HThYgHzO0s67CYFPWGE+bHU4pvKc1VyM0Znfyhp2FF+LqN/r2UGlJu38Pkc
PBwNrLUYGwvwcNo3YLrK61ZCd/0C3uhGDLPqTZR/5d/DtgWcRalUatpw62JmktCw
8lRjJ/o02c0EMCjoMxUkwW1rXLuxiAET550uUngC1mAkNEZVYSKJDIbfqbabcPwW
FsmIDGw9Yd0q0O2lI+XYn6sTiMk2cYUMGlRp9xTh4ikrTR//9VmvCGHjqRjNksiR
J3H5jZHf31/fyPu4Fv7XmklLu/mSIpMG9uHv4+rEwQQjtvyNMnWohI/iMTmkD6rF
31LaCpWhw/vFNsyXIu6p9pXdrUc99ElBct6t+uDTc76xj9igR7M5+5vrRWCbU109
fmmMoeQcMpuLHouT8Zan+05Us3Qmm2kak7djt4xUXeacbAGGY3BnnQaaEi+9tZCv
0M/CvyBbHNS4zWB/UWXGjRZyJgoM+h5IaZaIedQ098a9hYkr2DNJ6iT0tzwG/uZ1
3AmLLxqraG0rBifeXDXL27MQog1bltOBLRrNZZS75mrg3GJ+VBvNZ3SlkrUWzIoS
qDVHEWI1jfbLCj4fsoAmM0DJBTob6CY7Lo6kEEbEfKh/EZ9BEsEe81khGjp0XLDs
nA4fePkPRFRcXcc45a0a5UTiRZQ4APxTKFD2iG0pryOw5OPe5Wio1DcGFK4IS7fP
Ex5FzB9tx5v3YL4l0v9JBCFEqkzXmEJgeh3xvhC3CfzPx8DEiDspBYUPSxyXCwK/
5oWMwAxwcMLUBla+pbppg6q4Jlnn7NeVLRM264EcnreVAMlv54iYozgmYpsxRRiC
BTFDk8nGjhf0OzxHIVNv5K4zrAGMXm5cLUO7Kn3vfGOXcPbNtxnbtSxxkJrkWz2T
QymTZY0sxH0p5vLtgTZDolKs4LN+UNhvkNGFjNobSaKjIiLSvuuCYJEjMyeArxQu
6no49sotDqlZk74gsDyAtkykaNt47SHKM+THMGLiXsTpgixh7bfqQbm4JDL6nEYI
AFMntUJxGPjcyhNGty0UDT/H2tFW5/Aynk17Y3SKyn0JjJqd6aX+3s8AcSU9eGl7
jVSCO8zx6QNYka4Xlmi40jnBNZByqLGLMCTXiL+HV+FM016EFaDKQpC0N/sR7+sM
OTJKiAqUGtWC3ZGGWSgD14ei8qcNq9HPh9o24/acVAR4j3f7XUBQsSqTIGKeDEhU
aC6uGCkNM4u35OJYNFrATQ6LP9JOpszTHiIK5TfUprB1Aw5K5pu179We8SHn/aUA
kAbChFqSiKWBVMS+dODBNpBwR9LsTKGm6iS16DD6R1bFWVjcl4FVAzlmLDafdsPS
zm9Qrz31WCb/jHPseSTt08UczYXyd3APkH3VUGE+OOrfwIEwA2zGr0ABzlb3MlLJ
t1evA2nbcH9H9AqSenzqlieXkCW6RMk7081FG+VDP8zga+Qsnv7tuAPqiuk9Ctq9
87Jk3Gq7K4PKHBJjDERvIP13rXloE4LezA7Z93B3QaNlfC24TxdjUtfnGzxTJ0tU
5LSWkgX48t1dqh/q6PXGmu5IxcO5/bw+fSzulqzCtgy/ocAroNt5T2h4aF+KEvT6
3bsy+tRRNzNaR5S55sHWGpp23J20TpcWEvszFemofpjXivbzTvsDgi6IlZvp7e2l
v7/4Z+yq5jcNi8SSbxhBJu9yeYacfK+u9jBaWaql3AegnzJKc/5xTIh80xi/XEUP
q/z8u7G5v3q02CxPHzcR2KV2QwP7GBSTxdDf7qMEr8LnJf/UECC1TAb39m6wOwQ1
NKoqWh+QZFOiVmpad6hRt0IhKVWrSP1qWcvrCpIaf6bxetW/DwWpyq14b03Ktrkl
cMi6L2lULiV8T0j52lXJ/0NJWmqLnIIUrRphvG17YziGVdcqBoj4VO2PWSR6q+eM
OwAFQ3pZqCjDEdQq9uOCh5O7Eu5Fys5lvSJ0qa5atR0rLLqJqcv4YouIcEWcxPn5
vEVtshQvFWCgCj3HCqle8QRlAkYHiGpVdY+uOQ1CHW4jziXe0DSDrQC1t4AlJwTQ
bot0DzXa0LlW3aZfDbUqlifVh+aJIl0iYXO5ylTgbP4DXyN0EmLIA2d1ONCPXzkF
ntu50P4yt8+iiCPxYP07ARRMuG85ihdwi2vUrZUlPsdKvxyYdaiMzJMCicbkw02h
n1Sk1M6amRkaKZD5vzNXYQuhot1BcnHHqXHgzx637GfoivE4qnYDJxsa6v2waaiY
Us45oaYRRrkgSYDCpht3ShVSqAyPKI2WN9+TK7XDQunHG3SFT6Am6y0ojAoejc+/
TudzFlkAc+ByiEos8ernyWEu5iqSbKeiYa6cBO0DuxlIpE+RxNkMgp2JCRnshKuk
RFyVSEdtI9ek7IkPVbOgRC7UOzGp9/IynfJcRQ5IFSz4FF1kUTYGroqWQBAwPdZ2
wC4A51JJp29J5+agouEen4pUoZeIw76V46qtiwxyxPMNc2Coa0zP+ekgBMAoJ+9S
MHmXhpDtLKlGI2NhYVPkpD1QCmWgKYYeKEWjEBs7msEjO6DxDrdXKpf+b5yMH4gR
Pn9EeaeJoR5ZGqcKNJXBWwhLWjV9yThb/Ffu35p8CbRjGe3qFiwRLFJLeemvshuV
ct2hLmXVtOXJsXeS2TNx7XSwwGR3gK6dqhCJ8VgfLOQgzVAacbNO5XOXDZvw8RqH
TtqXVngeR9AjJs/taM5UJG+4szu6zRofISCGH58Nj/RWrpJzphFVGIc1eYjaX55F
EttTmAu+E4KtADO6s0pZOba1NySNHlD/H4vz+tRxWG/+T5J8qcNAOOjR3AY3uLDP
kzI6gmF6Go2pFmnk/UCKYvH+96ay6Mll5olBAaKzv2qU6knOJQTXkER9poW/AgtZ
sINB1Y/fmMTtTcxj1O4IDGBNA2H2S6mDq4dg2Vr641mT4UCIsQguJKXPs2DKllgE
VmY27XCDuAkSnNxoIqrCxgYEXSC/Ri+obRY5k5dFI+PqkcDJIcp6Nq5ofNMnU9eH
XvDhELuTehhunks+0mwbsiwZ1JiNjTS/W8lQaScYqBXwEv3qhGttjAkOBJZDFG/Z
mhSKXegad11gl3HdoneHk31Z1630J+TsKAwdI6ZXdN9u5dXPW5VBWFvA8gW0hrLK
k45ElcrYqmV2P7Vh/fFONxplmMA9LPR2CUMNbpqfRMLJBf76+IosUy5bpzhjSgzu
LzeCgZp/iTWz7lFoyqGM7JtUBzFVK9YLmeaYQYVxY4fjtS8S2flNHEeyAN6wSTbB
COEgtNY+c3PQjgj3jgup48JwNo9nHFL7AKlaubAM8j6/K+L4zi1A6zLGtm6/FHvx
c9kKQtU78fLyHAb2oCU05Y6Ck6G/HmLW1fEYekotYVdBQLfmWHXHwhVRja5MiOs6
Lx2ohbieKXMPjrG7AgsNjT1Jxs0dq17hdT0P0LgTvDvzsTn8eC6MgLKI5SIWfB8T
6XmUq+FSjeNpNYpdLmUEccIiB46JqIPmhYoBuKDLU7QkakP5DWfI0cTLDKcOdgLP
Emu7MKb8iAfqh+Xk7Q4CVWuckv/5bRHegTB2qVewIYb1Yr5hI0L2IJKqv3Ox25cW
L6U5hkKnpsKMLo0uots0f5bG0NOvPSUFYXZzZVf39qV/UaFbP8SSa6cZHUcLDwAk
c/KQoFEYrVkFtg6275whYWwDrn2EeAshECehreaddH1VBrs+wTJROTAHeENC1reb
+psV/cQb9WRO7qSLes1KgFTaWT5oOaY0PhMG+XECgp6oUBqcCdDutB53qwPCnElu
Y5N/h/UU8OymeGXbg9zdf5y9AYLTKaDF4mlPa1mBmNr37ddIeOKuXY3983/XcuCS
FuCPEjl1PhWtDJV5qt1UmqkOp0q3FaDJi17uiv3BcVQPyGshtNsWmX5cc85eaeO9
uBfVRK8FzGUUEGM8CkUqSkZe57xlsiq9LH+3GnlcghgjbFnRoion4lfYrIvVJXQv
z3li/Z9gprpgWUmXw3E1MzsP0Dk35RuvxE4xDV6HfL4jbS0k2K06A4rvm1R0B2en
7SjCKF6z1i4tBTO/585+isatLuGiu00kWPd2j2twvn+qq/u0cCxkkLsgO9JBz9+3
c1noYF3sN8/1wYkWGI7sMUa81qPleFO0N+FqfE/D/p7VOU3AZr5Lkcev8XAxqiTW
GfT0pHzDy+1sK5wwrlHr69Q+rGsI8npx67tKWseaKXes8CNVJBkuPXkDwVgC3LER
x/NHjfkuOd6COl5C/wyBDhbAXcLfmwwqV2ONFb3KfiktQAZceUp+eKahnfc6QRx2
kki99Hx5zolNechqZDBfV+Fb4SvQYPsabqJB5eBqtd5P56hsGzTgfeCWoQ0LamBV
5FKEAZ67xMSQwbpt8nhScGiqMO/CJ5e9i/nOPpGoMkvV4Z0mrPX3BxRXM2Idoxxv
PucRubeywJeZJq6fpiIV0wT5xe4WRXbzAq6smR0vsyce/3s5OhJRZcqw9oJ8MXIZ
54czfQGSyMMbTHLq3ix3wAqU+RVwKmQVknn1qaUljF/P//U8Sb1VTNahYThFLi10
m41tbFf3r1sLcDILounxyn6qXWGBDr3PoQ5r1pLaxacya35g/ljrj38kJMXquenk
PDcjA959VW0vIFP+s0DAaiRS5FnqcvSu93Kavr5rm9HP/NJu6XHd9Xv2IjCZYh47
6gQccRIup97MIZlL7RBtdHskHlI7tehFhZItpNUvcKOmUu6fKZBRhUML8kryeGVV
IkOX+wrlOseWNEZ5DUf29ckwKvb5M+Q0PpwuSRKCI0PqPUctVMPRaNlvlXck6oPQ
Wzjf8t2yyRtJuowA4qFbHX4aShRF/ki5BF71b0l6p0NvTfgDByp0mxrDBN73H63O
d6J1hXa2GklQWRvotmQ3pOpsrWIMfT+xXIAz51OhXfAtqa1ySHjz3KzMzTfUYzm8
518eTs60SP3Y0HaREJx1FjCp1B6e4jD8anaeI6ibMl949UQ7pOaC7rcvulBh/Fjq
MAL25M0vuqi4OCAJOakLlaPQzMsd6JTsaQhdqthaWh5chaB8iT/H9wnylkoAXZrq
95v4Xz74BDMCMUEWfcX4krrHZp+gSwkq5l+M7toYYZg0gzMrCSjMicIoHhALn+ZY
oX50/nCooFwzH9V63tpeuZePzlRrXsBYIyI/9dWYgaarAoCzTgYzCRJ8Alv7Eonc
5l3Dw1qqgfbzdc375eksgNxS02IjNpGLItWjYgqBS4p6IcjhD+bHHd5A3zBwJYTc
oyJWp1WWoLPjUYLoyj4qxS+GcUiVzJFi4Gmrm+pszpDx9Y4/frLSEiZZdZzn+8yS
RcD9rM/2kgOtkqWn7Ik/KYGdJ4/6xsxQkLh57Aqxg0pVyB+xkv7NyDZqQbGwFimn
1lMjIiKD1D0KqAYMVfbrOwH4y2faKqZFAW2xJk5XzmLGSXz/CjHErWO+wbr129b5
phYQpZrLm5u36gaAF7z7Zk7QntoBwMoxGATYzkBGjUXnpQljbfd81pb5RhPteXwE
GdGEaX16FbDYr32gNyyxQ2WUGtMTgvXSF1Ril5bFr3zIou/NDhNY9ug4u+MkvaO7
RDkwLC+ER567UbUFf0/SjIuPX79XsRVSuXYdt1tS+SK2EkmZbr/Dgja9EynWvHwU
o+BVTLYGzCpwWX85Db+SgLMEQkebU9aNV2nf7Qcv6ibgX08ny5VGHMMUseBVYDBS
WTzC2TqYvMcvhtx7FrFIUVVAEoLD1urw9ZTZ+kQuuBlux9vgC/HamZnhDTOT1jLg
RXomgCswzKw0fTQFm4CphTQ2t0wgzWO/Jr6gab/cu9cbECpc9IKTST12ajTLDy95
qBacDskN92T9LPC/yHWntani4EoywMRVJ3jYnwMKEMHLqwUHnsPHKRvtGhgdSpZP
UVAytWXOjZGWpDuwjyyWFHWFIGYPEo3nEhIWiwUf8Ah5ehQCezl/fq01Y81ALNTT
XFUtsqisIP3GShjznurj0KpfsRjhvWFAHfoAkFyfwzToRhum1IuHn55apCGc/jeu
8XQ9o1aOPYtrH9eh+MLdd89TAfXumYLUL4xOPMUTiIpWPqrF81VZ+MjyG21exPWG
3oGlPwexnsVNqZAcWqqGp8UAp7pR6X/pvVOPJ6a63M7Bl0z/D6WzeMtgGoaNQUBw
/1Ul475xMFU9slSXT3WAi9yxLAyzwhgDesIq7G+naUMydab60R7IDZTiWR5MVB6a
R79R/KSD9gfJCVIl5gXcl/M59EO0SzJ9PrrtNKkE8ucI3nUgtGbTcePEJHctjpip
R55I0OMdlq3+Vi4hyutkTb/CjHlvm8oQmPkCm+q6oZ0I2bF7HPSgSqXN3lxeMvgP
1Nyi1u4fOj4Kjg6mCBQWUm2C3bk+55ourz8nRJ0qYQLbodorqKqIy1/r84sYvCn6
M+7v9/PSPj/4fCnH7/yk8IVE3XusO3sExDrjl3Q4ZOhR6dMLzhy69d5zENPwgLl8
m+L5gx5W7LA5f+49r6iR8GbpFrxPiA1Uygq6x5c3R3z7q2DPebfKj89BO/lVVPl7
6m+wDYyrq3liSwDpD28q//ksNAXNhaFt55tLV+E4DCcy3DTpcNa3lkw+nNIN3EZj
uml0omE/FpDW4yJkyUAqsMDxRV4+zVzDmF/hF8BrcQDiVbI+ikJgTaRt0xR0/rmd
j9vikAciYjUKpCt/1bzP8CsGR4wjQ/VrufXJpkVzmaDFeLkg2RhWn8D1Nii3XqyK
RckVb6WzZsQP6/AT4CTwYybhBkl3LyaXjtiffVxL4JtOgHDSkUfKTFWaWvfNyZPi
9zc+rCDENwrCynSV+roDcATM2uvZvPnV1TiH0igTTHu2SWYnSeOqrLpKdNwdmYpP
aX6OCHDXV8QlvhcRLSxLzhCa6D44LZTL6i0W4QzX18WoYEGfuA405c7f0aIHC+Nf
a1bvLn2olQ0j+bFv3vQa2szYIngX5wZNu5DpSN5DjKACUgRUHYY7bjUpVmNcslFb
xPV06DjGV4Its9OTFj2FZ1rAXiH3jjb2WMn/OE64JwCDkLQCb3miwxSeeHM/iKaI
wjHnN2oKOEdsxVyRRr9aVd2yPDmckdHwad7PXLaTMOmRQx+qIy3H5crkJLDyDh+I
YhyQQzETnjPvopcYmkNT7eU1rz3+UdvkbfQvsuYDIC6oUZT1hX574XZy7wGM6Ghy
8QfJ18WHb0KFfrf7PT9C/hIB9XIpywcWLWjslOgcfnaD9NYcE9KFFIYRwoYCsfLr
WJNkK3hIjFj+xQ/Fd/kzCzwn5Mytgxb+VES+beh+UBjSZ/f7VHnnI2O/wbVrGWM9
pYKF9xe7eRiNw34tI7hTmweO6Q61wHPq7C8bynrujhSKTBSx7T3+PX98KZJYvG5A
QxPbi5aT8YxCf1aPDDaWmK9wzkAugko1UrmqvGvMOerg1jbgRfStw1Sm2d2nYTUP
06xwO8PFpdFei3T3aXaGok8KFKf7VP3mu+gMCxuGax6vuLwhFylH7iFnTjrtEjN5
xE01hxQpHyVsnab95cy3OHWPB+7eZYAPgAwf391iQq12e/DbaD+poHgm7gF/UU+s
KsQ55SNgD/xJSPfPMu9FfmqUh0c192KR0uXEmrksE+qkbDpEpy7JUzqaNNoa2dVq
hIYHb46ORQ+5aC98DdIRuq0NhT5/9a91GBZ2dPDSl8n8Rl4sWOaMxTF9pmPPMMl1
FhPH1ansu6qIZj380abkSHNOv7YD/jVqzVfpSAClLx4Xvv0AQu1kwxmipVZ9n62d
ZY8eZVgbYcwI1ltoxlMqLCHVh/mCA1sP+rqr6W1jH7vNIj5B41XLlleIYM4e31uA
KHs9VHDsOfur25pEE9iM3zXPhPU2Iatr6rOVWnQOhxbSJKOnH7NC8SrKE/0nY+4Z
19Wu+VZCQnDZ7CA+SNpOghQE9gv7bLGctd6jGsfgp2vFOqiakxGOsll5HCbrMig/
VGDM3JMZsbOQsSujE1wdpBb7ZTzpuHCA5RHhEbDAyzbt5C6OJaqeLH1Y6yBCXC0M
LQaIZJ1P3GoIkU14nmSnaawJ48CDEq8mt06LGA6yFVxilfuwL2avF5biMjBfZ1jy
JlykjsS4REItbC/T3mHC76Qz38VWMr9enV04gEsj3xxR4AeRHdyNhvH4cEcmezZO
y4pNoB+ENG52K8v0mHFLSnwV34TMiTXk4Y57f+Z9+hPDbemKKUOpNNeLr+zVJi2z
NerzYEmqLlFSvk894mzrPfsCtuGVuMnJgib8IUVu8VBY9wGIH8XWPlGiAnqkbEkX
eamPpvBCNv5veUQ/8vh8RqqR1AQcm0k03o+0ooc3cHW1iRu9dDonzaMBuTpiuia8
Isx9K7PvEIjByaB1uT3RbIPJAs9oAlDF0e6WU4on+9J20/eUHfwubhU9EEVELpBV
0mVlB8uHN7EbisQls5xd9ybQPj1Az3JS+3s7cX/ib+U6aC7kdR3IPKej+HguVLPC
W611NQee7Y4D4pu1TRc8/r5HObWqlN26FFzK13sMVWMjgtT374M2DveWy/QAln4f
KbRJ0j5j7mGqKMeqizFmsJFe/sVD5BzOq4UHeb+H3BmlCjo8MQ5y2kqU4A7B4Z+u
pRJIlI5GQpvsRQL7nIJ2iHdTCZFU/hsFb2ZawzCMlcGj2wa+bT/++95pfKyXrVq/
Cb3YTq8Y6xMnA7qPwM5bnndHLeXEFNW2+JnR0/o4tm5iNLYPC6iZ8Zg6bhRYwptk
aUVODmOAKyQdJwVjds4sYyqdxFZj7zSeAxPxgUUXzl3aqStgnNpPgUQ9zNKTklPN
6V3IGHCyUprHTw3xh1MDgbeZBrV5EUy90vZTUBGPPnsUmDezVM2vQkGJd9XYEZHP
1i9ggOVMyudb+ngwA8fS1PXDLcE0entW+U7ynkLFg+67VoyQ3vOkLoGgwiJLtMp2
M17dDqx5pPuC4SP4wJfHMnxlHslUw5xTKB+n8XdD//qs70ydlvcwVKRC0gXiLl17
KRCPbH5b9bW40iziXFZ42iCFU8uBmp4TcPQ29O/5yJ+az8ltJMMj9mZrLSscXUgC
X8R9DTGa+Sj52fPK3RONeaPzwOmCx9BvqKhA0fSaLrQZzk+Ht1zKMhGj72D5TFij
72PxJYWf95ao/f3Hx86RhPW6yXjihSu1ATyIjGmJPplV8tIU+9/qsykcpZ9TPNvt
PvhdinnAreBGpe7DWeMk8uU+8eB/c8U2qgcBFjvs/F6Qcl4a9kQ6JpWaybkiP9kg
7P4isLwe9l6r2rGoMtKb7MkNMGds4J9oaRXWgy88t2/atw9knXiCg37qIZnnbIEM
gnv8qHq+iQJV6gCheHSBxRpQddnETy99r0f8aUpKRJJO+OJKMBN7XVQ8RzADioXQ
oYGExGHKV+4/5djKPogGMKfVYUnpRyV4QXa50VID4r8y7e4VUayc3nbyy7ZI6fuK
kEJ4s49b99FSAbKOpuSZOqFnotUkOjoP0H+KGsoxE1EegrPCuqzcqC5QcI3N6BFA
kYP8P3RVACtjrY8O5rdwxWzwRx+Bh9Lxy6bCuvYETHGq2OQ4q9jlonIGm68bBbAP
pqxYmeXqG+PQ3VeabM9JMG3dd/L8+za+jzPGlh1WFKuvim5xwGZ2v+qmwOjASbSf
WT/DNoJBD531hhzvpjj3mjhup70E/Od2L8WDGMF/fHtqi5uslw1uAGE+ySq2nXVK
BqiGHjF7BcokRCRoXdPvyGahR/hSNOgd/3QcOZkXCn+k/rjJLsUrekN5wEDGsaeg
K9D3DYxcr67VO4kdqqg4HGZjwFJsmltz0/RnZIw+JUOmHKp+1a1rAhbaJ41FWAXt
4aHCuRFurVy9L11JpzwXsK+9SQRWMLCitZdi0RnYE31kcLhI3xQNGNYb9IAfTU63
Gh+KTMCwryoStB4Ewex8R2dGRrNLb1HYv7Yt2yW5nfPQ8S4qbGkFk+SFgYqmxhmT
UAaEz2/JbYBUmJbz3hEJUbwibhDINUzfb97kIPV2rWDzmTkrAwG2zZm2XFVYbAWs
U7BYZ605+cYyF7upGHgM3sxxwyp5PpIYBbPr2PgwAjzlmAkxrWHyFjXDGMagJe/A
PjQ/jkFe7YaykD7pyJHgk6io/vQzU+SVyQ+mnKIwK5xKPO311WR5SFwyojJMZZ+3
+PY3eoJ8Lq/vz3dzCoPelB2eLxOes/h/My5O/pDh0qtcpbtNJtTrJeSvvNET+vzw
ku8ZTbEwTeyPg3guP8WlMbKcWgg0u0bHHmrn4t3bFSb8gF3hzUpW6aKOQ2UJ7rBV
305f3pNvnKTT7Y6Xd41cOISZzor/lweAUvHUQm1exGqh/QhU5WMvK33zHM3z3DWd
PRAn8peLbHbPgb6XaecHAH7K5B/Y3cruPu2ozOPFD1E0cyUQJTCnmUgZt18b8uE7
SsdkBHdMrAbkrlSR2rHhxccvMIoQ1fj584iHuHOi2zHF5rfpeD1eaz0WXNfBSerX
70OnGxvLKlWWThzC5QXlnFeLI/D59/nNGIExj9yHB/+MAfnZFvKT235J9raH6Z/6
ZpcPkXawUHZGieereucNTC3cjmJRZX3ClTmnthwCRY5cXZxi17Gxvjs0PJ3KbWe/
GXq+7snvKVKOh0MTsDtN9Ci1qf6/M+Xu9CQCOa7ifUws5jTxsc+uGaGyu9Ri3nwv
Y8vk8yJ0wkG26zbwG+sMUaNnIjuDfdGfZna+mjtTqbtJurAXm4XFe7x8cKs3SfnS
3V/exycwHvxCYRkYlntAc8R49GvjApfSiIyhcIU3EbK7RnqIY7KArXMqzEIVUyDT
B87YUq9+gsGNyRkXidxgzeyTrEwHuenb5RvdTm0whRH1yGEE3HSaPUPwKRL1iFJF
sA46sTyH/0sC2Tu8pZPOUR3jo01XxsrKI06RPPmU4T9pDsDM2yOFALpNC4ADamFy
2J/Kg3PeC4Im8JtPLbEMPIDcElTYDVDVF8JM6XvBHu3L6VYS/j2b+mrM5Q1XgOfm
A+3ccBjNzcC0xhN6vXFdD5+J09Fy/o7w+2JPPm9p4xHnoq6/8pi/dyWzYbSRCdk9
l6WX8gSS+shgfBH4D3I7QXg0VPq04rWee/1+keTlAYWyGj1ELI9rOv8kBQTT9g+j
ySz4mrlDUCHBcees4oi8M3r+nCck33xlAmOKr5WRKgY=
`pragma protect end_protected
