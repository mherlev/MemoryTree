// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:52 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
WGYrUwSS86qISzPnujz00K0GuhIoVjeVZ+rhLGQ1SwNjAiHpCs2z/J4nFTUvkJdG
KsyPcSKn8DrxxO/mXMXGM4Uvsr+zFo36psLlCFhDrqNRYdIfX3kAeROHjTQDbhlp
UH+Iib0b/KJDdPXWXPhvjyBmBucvIUsI6WoEq7fbWkU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5424)
9MpdG3v0qmg0vcrXFglOJeSb9GM2OhujllNz8thQNJ6Xfp60tWohi613hqyFULAq
ynYafCW8iKzYH0jFLnbiU9WcPRnhknIT2dc5/m7xM5s4gWwNlfAzhaA3OpibWktJ
WeP/AKIQjeCVluE6Zm1+hyWEmGydyaSaiYQl4hTtDH45zSoIGrVfHjYP2D+pAlL3
IzcVo1oBQLLTTkVxmxYFrf0qKtCgseaST9+wnXaIoeK0pUr48vZtrKoYEMAkG5NR
km/E0t4zxhD/5QoRcgpkVxQDEqAsAJVdw2/EeduYWxbbtPdOQNq/g9yJ4lYx7/1U
7GYsdnH0eEHmlI0XV3FPKQv0o1+u3Tsn50ts0H9e278ZvxeUTqFTitvlyype6rbr
rpU4GBirr1oasS395W1Xnx720yWy+4oFM64jykYHq+9Q/sK+r+YEdZhB3dBdJveG
sQKeipR6q/ddtnnpJvmQO0d1KiJfK6sWqQ4fvPS23iKRnaE886F7uF9r4LlsXsK/
fgtxxQfNgtMO3UnzOpxC2sxcUXOMwMkUMK66Q/MlF3jLYmRZB9r1+3sWWwFFrisi
TVRqQdG1n8FszRu4SM2QrYUrmviuKkFdnnFyQbaqfzqZ1dC+sadLB8ueWYFFw6oq
s7FKMrvaa+33mxPP2/td6z5Vm/Hsy3j5cV8ZODXpYOZw7lRaHwpqUECQbz/kXSni
MxZkx9z3XbqE8fSX1isNmW1ntEQGa3caw4AlNrfBPGFEMAb/SeBpEfYuNyB4bDRC
MJsGvnZHSSOabP8H0tnqQyOWZNVDmpXD56Mbx/Sp85lrN2UsItGL+ySgES0+bvmg
S7tWzaf7wEDMVKtFOMW2fqWtoLmZkmT8mfSrr5a50D47Vj/I/hOmXEvb7crEYrBl
XYH6kWgniLE5DdankrafNMMdfBQbiYHmWQ2YgkxqMrDbanAWnMxCKK187XiQpXGG
DChL7Q/vN12uE0yg5wBmMbvWYxC/YLmUn4HihBUwu7UGeRtGvHhE+iw/thdBgRpB
xVKcsKPgzo6N4R8Ep3y5dMslZWELiXD1frZfLz/Y68hu7g/jmAniFN7wDIi2LmVa
YGHJOyGApG3lqtaFKMD9QL9e+lf8uwzr016tJFYfGf0WQPPievYufoGBEi9vxrSy
2qL+qhrqaXekC0/EiPLo+VnPmQZa+DAmSVk0Vc3yiV6EXpogd5JBrjEVzea07tHe
Ft4tE7GXHJc/acR2+6pULqN1SulbYT3XksCQhXOKbGVdZz3AZN552xK4NRzPbYFN
nk1v6B/QumsL09836nldUK2zXn4d6KtAAIT02ecnUXBzzbh9NqyjzNy0SCmhh0Xm
smLYSfjwdvSfAa9R6CGCw4i4UC348pc1xUEh34Jk4hYNW+Pa6sJ3Vo9yz1nAdqs7
B8wAYAihHJfuYu48ucltuCagybXkAe3FNl+VOugBFRaDponIitJ+FOX1J5Ld0274
jrMyIx0BmRgUwBMCbVz0uwetjskhTq0xW1tZY/PeGGN1C8LKgtTlepMvI/NnSJXj
GrtcWEQhRqUhCwYgYZpG4EM6RVjH+KUHbKtHH13HihfEKTWyi2VNwl166ESCtjnm
QLCpdDi5FfzoxbLhWqvhGkIdkhWNH0P+2BJR6+ZTGcbpxDHBwjDc54Jof0KLxSnh
874aQWQgpiyOfq9nxJ4q4rLyfoLe66629E5M7JNGpQYk14AMWmSzpM+VCFXWJXAY
uN9GYD5FVrPP1Dsbd60Fkv5lUGM8fu/dRNulO6gd0vT2m5ej8a0TsN32wxRTyGDC
08hHA3HuJOja+6+nUuquR7NOiCsPXAV3+OG+MwLHJ56sAO/IzcVW5r93leePX34N
lECit1zQdB3qBtdbAgrbFbZ0QsH7O4H1Otsckhl4STla7B/ia4xOeyUDOKz42PfQ
PdTH60eFguF5Ha3sahfEMmOgBRbPeVlUbf9PsFFinxVdpx1MtS+TF++c6TB3bjTy
+vVtgXXlHOmvydclyBk028tz8epnQ1uIqzFAV+yP42+bdKRfE6WGPNscICbiHWF7
svGDHEEfeSJbUPl8nl1NRh0rTIHDqc7bi0TNGq53lfCRfO01o8UM0MuI8WF1s0Hj
QNopg+1TMvlO5M0PgzpMdi7iuE9k4li2sBwZIt4Uu8GlrbMaChqTarzT81IvYkT4
hqIGNW5TNG+lenCVQxZy0a3rtgkwsz3rnLfNuePvK/PuyZX/IuyYMthCoskkgkfP
xCZC5iXLz9/YWx11kJ2oN2tJEaFi5HiOdG5HQq3MwXekaFu8auIt41y4oWpbctQU
Nqsq7nrevXwhI4b+ehFCVOaua8xMcFLNBSGGccOPLQZYOEB3QBvFB5yRE7EXHWzD
B07Fh7/5tgGeWJguKRU2OS+SM+UYed0+e8NlksWoeNqXNpZKqoBoRKbBj+hVrM4S
R4uJxpkalPqPcUZXUBkybE4pDV7g5VtPhW1neMe47RLIiJ8uGAP4OwT7mbeGcfxa
g216G/8ZrS8ImAYGN2sxLu6kYc82wXjIBJLLB7OTAPIGpd4ufVYrtDX00F9lYFbe
+XOclI7deBn7LgnK74WQx0e/fP+MiizFMkd/TPk0T3n2d/ADO9b+dQ7dyZhyUMnq
yq9u3N+sc+J1JnIQtVWoa2r45OMq5yfOukIu3y65xROLt8WutbsgPrN1Hlv4tddh
szGne3ugG8mRFVoLltRDRB2OgC/VpRnIstn3qQ0IKYsRlOpaKBO46s6AuKwrS1z4
EeJiypcPezwNPDHgPJOD/zac4q5cJ0WH86A88BdBV0tFE9Dcx3uRc5aJ4gGgmwjq
KLtnvC+/HwtegrMZyzg4aGd9CmPxGO5sZ++i5HQY7zFirvWLYbZxnJGeTj/pfp3y
TR8f0y6qz5drNEdg35fory8+t+hYiPOxIFq2XbE3vVg0AW/8r16J+B4d4Dw0W3QP
8GSWeG1DCmK32YePcJeVWUIgqAcWXOUT4VJOxHiA32qDvhSIw3l0ljC0xBro10fL
MiNVSTSZRbfY+aSdEI8rcYVsnoK/lK/fmX/rKJC9j8THX4wq8NFNJWIDyigPuTYM
I8FbhP1eSgKyMOziXyXLglmoWV114nUQdJYsiMS1Oy79w4UNpuWHID0K+3yRXKuW
s0DO10BaDVHJ23jxRERvDWMyrfc4X79CETabhVQqBR4u1/3ygG3xNWVgD/YyWV3O
dMp3H61mLiQ6nvaYr7ELgEkVeFOKgTPKOtSmrEhhfXc0+2abeveh7ZxbcfDNChSd
CF/0P/0TX87ddmk9brbifk1SlbDvhhqrJNDoYVigiID/CbSG5MKiAmIj51j+dP6r
eQsG+ESgiSuicvFYRv8Mz7C9yM5iL+w5TVgrl5zoWsUy4EUNYKpcB1516fK0RQcz
1ENdpDmW+FeMdiqxguewISxPFt55uN49LBEU0JTXggUeOmIMXz3i7ouIapi9WF9I
WyaSbesKr+BNnwq9Uh+Slo24tycH9D2xRSiWQr1CVsTe1KjDBJ0oDn3PRVGddlX9
v+ZWBDeeLGw8Hlnyl5aV8NngAWCeAYw+u5WKN2VuFeYBQ5UQxIqGmYUsZb3+pMty
DxhRWVs8NspEJdclFi0ST+px/rdbO3xgEwez73qP/nSDR6f/daPJulwAziini4iH
AhhX4/kM+hU5Eda8Vql04OK/3JzJFeQLoTfpU5sbjAQzIcUCv/T04ZSVi0prXU7A
LQ0tC4QuPOrUFVr8Vvz1aehEDnyDxx1PtRamhnjuve5JqdGqZn2DpVa02QmxAh2N
fz7EzVe+T/w4HBHWLO/qDgyxshkGll2Acu/V6iu7SCQBQAxlue9wikLN26Jh1Ufh
Uq06a5Y56PGUUr/fwjX3e41B7CuBN2lmukWq9eDvN/illJNg7n3+2RWTMRd/BH+U
IDuJKh4JE6kclcOUiqtX9w/Mz1DX/mVyQVjVvWGawVbvjUHpN7InEPkud0iY3soB
/9Ejb21YVRK/YpG3pJOhuXJRKfjY9wTRYBnujoHlFG9ZfQSTZpA3uQ529WK489Tn
kobaxwc+GSw5dKcClI7G2XTp8gU/VtSUFoxmAIynEAzjkvYGKcljVvkWCrxiG8Ae
HI0U4FRjZTUTasLTN1R45TN+btKBvSzVNghDOAKm09yFevy1g8E68i+sgyJh97Mu
GIrcVeCdwAQq/BEhFm2M8YrJsncMb5rWESTeg46MCNgdnL3MFhFZBom6xgv0p1RG
3gjiAAkhQpu68k+/h6geB/L4wfRi79tuIwwuG4bujR/zFmY2Tf939eQxsLKQQIWB
rcNtGpsuFkBeFiPzbd+oHKDC0ZHpzBN2N78BuPBO6N/HeNqmnuefJOEX3wA8u6bt
HetahpRpfWBzWZg8qEfPZe+5lO3wW9jhtmM6rnS4LCI8+zIL+mJxUOAIFjfqnINX
I/ZtvxnVLP2uTyHev+0+CAeN+BuSNgW3UNBUe8ja4wqPygg+3PoRnnAjsYBbmTX0
UaOG1Yd1c9R70UqzzD6R6TvWpkRvYc1cqlMep3YJR2dbUVmwm7cpnNoRQlLzwT4g
YVNiH/ySXysqKRmrG8LNBGQ/QcPm0J41RYen2VsQA93iLQ/Z69i/bd+6ymU2PYJa
J/5nZjlNcb5n5VEA52Ytpo15A2TozkCi9oT73JnkY0I371uOQ7Rk/1TiSqz5fU4O
Ub+SRFFYVpxQBFef1sJaYCImay1PPqIpfg4i1bapoW+c0s6qpPyEk/kU2tQ8fpJG
Qd7/dT2ZlLNAbtMWlAe9ueqPxF8iwO8dSc2ZUYTNsvBam74X0pWDhPWryH/MUPWi
IDFSBiE+CJlFTLaHLP/2TJYGlgYReS2m87GMiV3zxb+P4f574Gy9DWIYwlhZXdo+
KM+iY/Zzyd2mt492aXRx0ug9U5thrVK25pipC5MUFPkzakx+GtCRoDlyPZYbSysf
wfCURu6Q4VYx8ZLy3Qw4eZZabN7E6DA5ORL71Ij/RB1qD5elZxWRFKgkcGvXy62U
E1CzN8pc6M3Yf5KEXgiBFKHnNedDaIr+bdLQwQcfCewUWMjm15Gjh7WLEvn/S89u
PzEgUgYWH6ZipBlSXkyKEMrU2YLu55XmH/B6Gg8t4OgzaHPs/9y4gWC+Y+28YAZE
ZOfhwN0e7uwPoilX8BHjQYZOnLtigUobDBSrm2F7zyTGHZJ+OM9ofUe7qGriiFng
X4sqKy+0uQl2GA9hUKKIopOn/XPjJ6/iN00M4p6A246QaS+YWahg6/50aqL8wBfe
XmPnUsnj0WNLa4EpZjAvK+QGshkQ4IL13hP7lNcYn73mFZyTtYzP8QDAnC4D8gvw
/LR/H2SdlHzde3cDBMslUtIL87PhMpWfVj70OOHpptxX0xJmeTd9Em8DKYEYZWo2
wp1T+yaeg6PeaJVOAX1chWkwkT+Aa4ZH2+Bfq0Axd4Y6cn/R/R82D9s2C1jpFXq/
Owhvl3limhvjFNzGq89xq+zfnWt0ZW35hrlspLM6P5B14wiZaYYKEk4E7XVlPths
pfBUdqskhXXzIi40v5yfcBIkUEjZWzpUzMHqm9EkYpCsfu0iden6QaLEFljERbUw
qNVCcAmeWfGOMDJigdl+cFzFdnYZJkmTyuZdfCZc5RfrYvvLTD1hkr/vNz1N5lCV
74+1cMSn9AmsyY5z5oH0+mF73rDQqnrMBV1WnVMA5uMhr2eL7BeTCrFPR7IsOQDY
M45jxx9gVgSwYXFphmGYTqkd1PXqS69lKeA+SwVgklaHtraX4fkkECwuzIzwod37
Ar6RwDzUogym8QyfCnKWnydC0Cns0hhGgmbruL1h27i1NdW4QWZfG2d7AOjQ2WSK
YlypmOhQa+6UiXPdF34kRxDmPno69rA5dnknNG9l9C4CbkRtDryeg+mkkldlBU/b
evM2bATMk62Wgbt1RjQF5vhNkzfR3gkdY/cLyHLmCBJKIyJRtuxTehf+aIUFOfx/
z6Nh5bxbxDO0Sg4JtAgLM9CQXTmHYydrbq34DEN7L+/ZI3q4+K7BH3lHWvvbPDBt
QYKfxb4X9vdH972ie9W9jPska6P10eh6CHsgZmNpGLwENhyaaX/joZG0+kAWPAZ7
w4U93PTFJFskizl5eMKfjEJFFJevJ8ehhS/xR4Z2YRTtB5A9ndEkXr2J5q33AMmT
uv65BM04Uln8drv36C9l6hAvRVeOKSgc+dWX+doh2f9Z8OI51+6qtd3M9TDv051y
40TQ/N1CUYdom2zj3i9nw/6VpM5ROthVXseEyDe/HbQfJxiTmYru3uEUWqF/qLka
R9RecSLZbEeLdOekpMuQqMYLo0HKSD7w8OkAtSENp59ef5fh3rk2a+f80lt5UhvR
dggGNKEE2EjTC303wqOZYeFyNc8eoCWwSsn0UqUCkTRnFnnelTWsHwmR/xe+1e+M
3mVwN9CydCgiHpIKaNoLQwUD5PJ4tjYShjH1t+Ds+ycWQjCjyPhyDlH/MQjPH1iZ
Am3r11jpuRWwTEXlBNCQj1TTH2YfQiehElDb+WLUJ2bGAzQgzlR6KG64ll8/MF3A
mPcpEy5RwAlZh1TLOFyRUIuJLxPNfJYqKjgryWH3SsUfS/D6CvdaNNz4TrNe1JTT
OEdW5aD5NZt4zK2xcG4H/a6ntbKxIX8926GiqO3XPRb7afDRfd3f+uWOGYebXE+n
uOKsmsc7dPVL+xwOcB2siFzgwJzT0IQurmNN27mSnkPQM5F/EgBqrJpT36+Ky8H8
4C9zrQ5K/Xi4zSGUoPtyFQJJs84tNO0T3RDQ8WVO7Y742iePmBp1hIEu8eRPaa2U
Z/oTcbav0SsUYL1WRu43/+KbElt8q7jY2Fm9bu9dOKWMu2Ty/vbkErArwJoPSrAl
wrunXmhAZtqD9dgdysVJa82nhi7QFlaR2kITiwCiTvOM+NUC8fjpqTd8O8toePSj
JUHYznQrugis9VpQOKKcD1TGy2NXveWsqkfYZX3GaWH6bT2Vm2/NcQIjhqJfpP1q
bCcWAHQBWKa4JXXpp5R+zusAdIzdQp5JhvmMyBRCpc9WHsTI+X2TFkhOnue1vVfT
volRhr1M+ofwKCXEjq59UXGjf0fWfdV4QDZ2XaYxcoX7KyRLg69G/1iBlS8wqBSo
6fcaYzqZYielScD+DNMt9yzV0PwPfVr3BCTzSwqOZKi0IIedAK5ubMHV2E0ebhQs
TpIuMWIkS/Lwen2yFUSXxMqIrTdQdHN8aWA4W63y4riqfgoje7XY19guBDWC6W73
`pragma protect end_protected
