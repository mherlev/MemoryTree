// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:56 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
PrtvrKiQ1iwmVwej3BDaWVxOJMyQndq6+y4fazgy19M1O95nn+OtS0upjrjPIBDI
c/nT9z8LLCPeVxVxezSG4Hmj4MaImC+kP8p+q6uaPw5raI46AY4Ae3QZiPgFx6BU
hI7zIYdYfFYdGnfcQR32ODMQuddATm3+72e5074ezOg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5536)
rqZWnz6aa+KIvOAm7RDsCsul9fJTlOjcy/+SSLlJ6Pts6mWg1CLLjwUpoBrH97ZT
iG+1MD3pTDnwZlMvVtVlIdy8mxoGpav86zVhFyvA0JQocX0k1+zSfjXxOJpTWoUm
cEuGnic7LWfRsaCdqP0cW0Y23fz8Lyucj85R4wRBipB8OBZkNu5HX/NJ+xTg76Rd
QbHyZh7eaXha+kVH7+URY8xxQTC3WxKsyZgXCe2iywz597TXIjrsz70/xrwpnWuX
DfFlu3ifEc9W4BOk/YJFNbJedVH13BQX8OOjH8Ul1XNsT8y0NUCWCS1GADQgFsGN
tOE8ZlKlvAcdoNAo1XjDJq70Sk5ciPBGnmkKJljBFOKD1g+YM6Tu3Tdi2t9vmpS2
4HbrbxsenLoSITXWjlaQXlL+VXKq68+RBpVBemxbW7CBvJ+MIeOXwz+vYn+v03P7
6yn57KzZttre/ZaqAXj+VbynvvuHmKrq1lN6EmjSxbU7Jio5/EcPYtZ9x2DiQQia
JAvd7G9oggnYVZQcieS8tq6acyRV3rESciEyxpwXEHAkhj9/tKQxwuWhE0d+I4zM
bQUJ950GCGHdn61NmV8N7bWINbGcZgZttId/r1gHpiS26b/OafDE/YNEJwRdfnGR
BX7cHypgARk0ihd7bVfT4SU7foN7hxax8jPGKJNhyfqfH8bXiElaWJIyPSALRpyR
AWGOU3JY5PNZ3ydMeJDWdVf6bhn+LQWx/xFLgIiaZHZg+a+b7eNH+si5YbhIDcbM
hTyV6wtjrK6/fgerr9mpMwDM77kTlFViFZI/mT2B2DJNmRP8RfZlBLf+4h9+dZJT
NAVD7QYHdXC9C62MUH9F/BQVto3NK1FVk8ixvOcn0D9AXwrukHa2H4mREN1TS5Zw
Ahir0iH9patmRIbdri1SOOynURPH96yMDQrHJtDyAfwlrVbdZqpkaGIa3Nz6CAYy
qXRrOupGDBDgf0w0skEJCWjQkU0wK43xfy2mP/uF3HrcGoAMSm95ARwSAYShm/yb
CT11yajbait3Ri6SBpBk9uUtEGsK+FOrX/lCCzjf9UyhZVfguIVEj9X8ZwcpxO8s
/VOuOeq5emoEwcEAPdotRGSeQXj6hyfWENZRPa/shBQK2GO0iV1AI6qozl3DTKpy
T2UvHydqsM8ftsU2PB37b+PYUzGhLG75JhMcvuX0kXdsgY/+4x5IBL8wf7ei1VQm
TLH4koVetOfEf/HulWuYTKCKqs29Z3n8WymJQfBeOVftetcCZlmKYkIxf688xV2l
cXBpEt3/tDhCWNrLvPhAzQCPmIa0Rwo682UXUIL5UDSfpio/jmXUsQZjQxcsIIQZ
6SbEMTIHkcKpeXTQvQXM6rQHu2RYK0f7XgiIZbQnkBqw1GQLBpSFol0foBs39b8L
YS03ftPkE+CAo7eDXEoE+u45MtocHbpGj30XbB30ZUpj8kZvh327WipQdILX5fMm
4beKSfa7ex0/LA4m1PGzoIVOzpm4PKt7UmIjSoqGs8KsIHa62thM6yknRs78Ly5I
STAD3auqBNFMObeIAocKanYrhVXufIosGRtS+9oR7Y5Tgh8iGSOTekVRIOKQ+A67
1PxM/AwwBYzQLzi03iftjZl3LmTzjBUrHQq0J0zdmxCzHKbf8f9MeVkEdJz2LU50
iXfei0TC5ZPzZbnzZ6APYUYnJy+xM1ivNTP/eXRzxGvu31HWGHnbeFTIWSCZvdXf
8LwLx/wbILvRLOHOATSEkmXphcxdAv267DRgrLCxXNNBseyYFkXQBkWnXy2LodLx
MNxOWpO1R5OGhGkx/IXe3lJtJ1+kP8zf55Aa0y5kiN6lau8k+gDg4s9TVQMuvbfi
bbRlzd5KYmbeZ0xLlgzlV3atYHWzjhNJcg2KoODg6zwuPzp21eZNz//rvX9pgYeC
WAO9R1VfVgvVoHFwL6l78r/ITBY5eSnYiDRFjPFLsT418cK9Bm6Ah+Ic1UmMiz/U
y6WTNRctTYk2Gq6t3EdGgCM/UEVShPj3zuGTCemR4HVruEmY1AJ/N2R9F5U5AHCA
w3KKRODZwRaIqhQdg12RKsCAAO6ad74tOLtEK0B1fZ47lsbBvXHrNu02aJW/n8N8
gC5KV0grGB6Hi5aYhZD9w61fEhh+gyUxtsogE16EYgI/K7aqGvv6FcwGzJHbjhqm
JNARTdKsEKUEFnjcKsyvBq0bS+PRFgChDm0a0AOmBPUe18gyeqBXkhLa7hFRnyeI
92xwLdJwhj8S2rfXbi8pqcQXijDMy9FBfM9w/uuC3CcHwwNjl1hMRJCZhuDAGjOV
gqBST7lvYqNyFcSl57dqug1bCcUlwA2nXF98NbBf3xzSKylubGJhjaXr8Rjna+Bm
rRUBzZ6D1V2KJEDE4SVN1c3nXZnP+H9ZFKpTBa8dVOFRqgu0tR+RtzIlZH/Kt6iG
v1/V18WfYjx94lcCXdjDdw8K/eAWCExgh+sp7qUtp5xAJkgsO2ohXsRS3Yd7piBl
XUeN3xOBl6+jYZJh6BMMQHdsHhX/5TqwBTuAlX+dt5tc0Y1ui0QC0lfRcvvmR5kz
a6cgp97jyFHDseFsFSvh/7NZHA68mBK4AY4d1c6IDKUd17hvAQahkw9Yr6Ve6qM1
E5HWFaVjHwsAm6fin4o+t0CIci4FciCXGGEE8Pz3M4AM+iP2PYeYILoJMnM3ks2t
QsoG00HZ97jcgCbyj9H1066HzBxvpWyfnorC0tytfWz0STDRSwgI/87xqYQ4FDor
WnsSOx8stqULORoepYEpcbZKbCG9FtrZ9eiMdaWs8E2wwIXyO6hZezJNHhZvJcUc
uRP2RMHm1zysY4csJKoLKZ+ulq6Mal+Uvv/eWNUgiPfvRjHy7l5EX+twsCBSBccp
wcuTadKNlvlE6GRE5GRYWoVAQb0/aUwl2kAPwptFr6Qe/+SfJki0pWke2P/FOD4E
pj9agnoeLOt8bzS3qjA0MuYDs1TZWZZv8luLIPTv0YCeDyOCAZ8ZGaPl83D6Uf+W
pfT25qcEl65ordlwMWy10Xesg5+2dfCzi6zyqmt8v7qBmcbfu7f6kdKHD1axOuNd
4FwDRkC1yG4ntM2OtxgGrKrIoiTAIDc1xYPXuFV2CsomHsTUZj8mDlsskKaHinnX
9hGRH8NPikY2VmgqSjZAfoD6MKQzIeRcx02IjNsGbmVVpodN+AO6BacNbh6UGfAt
d0XmIzvC/6TkLnRfMBnzWtkb1cnL2RN84jBWknHV6Pr7iG1KzOqyiRWOTvHd+HkP
NGUWNC0uyVORavKAp0wO/LaI232XSxZDSAd9q79kXDJPwxolFI9pZZJVGax33Cnp
IMq1PDQIacBu4gGefgB3II5vagvxtOtqP/uawFJpMIXki3Kpmw5Qu72vbOBzJ5rc
JEg8oHCKCL/eMehVuNKhNJGJXHiSUGrZTRub/e1hvgGcdJpgoPEn02jplanJmN0R
byLyW1n7tVdru5W+jX3aSQgWJu2RytvlYYYj66CFLP2M/szZtf22UXsAI4uoyhG8
WDzHrU3AAXEO6UCvz5EVlKX4RD/ri+/nqxY52KOu3EwTgKYKUOrKF5dbqDYbPRfE
k1xkfenZ7diE1KhiCaa1hpvA2nYrFLVdM/1INoEUxTf0uGYqmkwS8PldgJiHSqEw
/uDmIOCrCFAbaPyN5lM8uEwBH9c4mPiJCRRAQlvMYYp9KQJzYzu8GCO1UnrGYZ54
z8FM48xfE2w5Mvl3a2j6v1SQolhHAQ7d2FIcIEXzWccHZv7Q+5PMbiZFVMfKou12
HiwvFifimswWRRKwLfrWI3+6kUWFHzYCMjd2V7GJBDPQsXeOyGjivu3forvaKFl/
XY3i0cyf3x2lOZptHYUzYfQ/UlYuGkpUsgZu1rhkyHiLVsRjVABgNOozgYBDINYa
mu2ir9eCj2xPnUuucePMdr0hqRap0ACUzEz6W0BQb3Q7E/Sv+b+KuW2X7wHn+Gam
KAqNlmoPL6oWyvMdK0vmnW9D53KfmnMPLZWKaP0dVOBpM/JzdQIyir57n/tEKWAG
FpuuBGhrpBoC+h1u/dq3wuije9I5+g5rxyxeJGTIlpk4H5kioU3N/Kqq4WHxglRZ
PYUNzcCvLY/eVZbyHML727AW6PombpI8DirEAy19hrdi9N4M6xscPefeVz3wB4xH
ZUP57gIPy8/Tuurzl6FCOgcn7QHa3yXyWNunh2fPqph4dxGv5u5tv/BoOKnGZbMl
1viuurvbqJ8UZUbrnoXiyLD5v+z/HDpBCWOqVN0vxEQ8ajUki606x9DtXKvP3nKP
Ynqi+oy4NObi4AU/5wcby3ClAk31AZLgllXOyICLC0Pdy3/YnIAfyP+PPB9468Bc
ntkkTi4Be1LRMuzAaL2SwQs8B33O9aI/D/H5+0YZX19j/T0o969/xh0j07uE0wkW
1gu+Bnamw+RPAl5XIs8KtLVSAGvD6qKWtLjfxWi5BBaZYB+Brj4BPMhW9uGoYolX
gzCGcl+zmEZJR/duJbaO+bK6iqvf3w+HF3Y9xFU71QsWzvZlE58vj2B4moJaHRX5
GsawioaggCdBUA0vqom/cxdTDllSEaZB88AgOE4IgQHAR1mBfxUqAXWruyTK5Aw5
75dSTyeQ96LQOibGBqAKD9zbxztAV8vfNpZARvnrE5KDCWDtoLYPl7L+AHSQgmcp
LAZqjy/lfUrycfIzoj8u7dNEsghePPp5C4RNfNcwZzRGBpLa6QTH1nqRLrIgu6cD
aFa3BtTP+MNHeJyGKAnH3N2q0iDZueNlsd6BhvZp2XGXyD/bso1IK/NmE928piz+
V/UnbqzdPw4ftvwOV47sjyFag+v4jkId2az/d+OtsC4ZJY78zQ5nUwpbR/1xWYpM
YpAFE2BhcemOYUuyUWkS64n1uF4bG/a/LOKWHQJ3AmN26QHmRQbGhexvDu+pC1+9
fyjn6irXmotUFb7ffajXH6EtClTUEc0e8Jf7J+uQtm9fmoDUBJ/LuSbYvD+QL+vm
l7q0aS7f8L9Oq8fiU1FYrJHcgZ5IMSgbaXJRTRf8mT0Jfm27iHtcWkLmQ5kBVol0
7cB+5XPEP2xjDEbw5+J9MXZ1TnhfaxYQmLSYOOZOO53wxVyg4gFonT7jLe6GI13E
VLwDADstsuE2rgEPRtVgnxBeE/jFmFPtcfP9+R73lKLbh+j32fp7Pt4ZW/hSS7SW
aA73D0PCBCpjxIKodaQ6rOGCEstUD1P1ye/k61s88W0upgv9INiPkebleJeCqv6L
m4BjMdQ0V9Be+KaDSJFEzpZhuOIZ4JRfBjiJ4G0jMzWQR/BZ3trdiaHHkoqajMZj
QKVufpP9MatSjb9VIeBhjLRFJxKBry/nNtClKB0+x9qnTfNthiEsbVoEqReopWRS
d0T2wJbQH1/lK9JAlDYYQi7SzNN+7g/NkEHAgUr4/3XiyeAWiu+mUkV3Gbvwzj5E
gboqI6BAXS8TeFPOrDJZLrA1JnUaL6zApwhZ7l5LhObA00dwdOsKESFtRSu9NGbs
fr6TXMnIXFaWFML235OL6hfpbCr+4B3z3OHP6TEtsqviyjweCwOwfQdPx/9zx/P9
ce6Fyvxrv38MyWlc3JzmTGIsIMbok26O/p1pH+/eLMOq4WGhSObjGfSEhnaxCana
fsrdoR4KU7a8BMa1NXoejSjj92BlUOb47y344Nwme0SyNsOiEXAE/lUZo7xSSHwo
X5mHXgv2cRxPZYSq6KOSNuX32IsDJhRkCFP41olzdCSaNrmR/CSUIZ6QUYwt2R1o
mZwL96+wyRWxMuNf/Nz9s5QJ25nXbAfuRnZHBXKwgNONxdkUO70dF3kASM29mHwX
6qcn3QokP23kh1KJugjaPsn9U4ZD99XfA9n+ACY14OZH8VxNeJi6c/sZqCpC1+Er
h0tDLOS3YUOv/ixSmGtmzfnC8kXxy699VP7j49+Tiv0gUmsONGRM70HrOvpXOloL
jgcuzzSWrkcMjG8NEXmNVZWnZEaoCa0JUWWKhgp9cqsRacGKtT1vdEBfMEMPOGWR
ThRSO9TvQDs2QJygAiQRuYglCQMOOQSBOF4fZq5GGT+YPRPWNWuk8wOC4sVJgXCK
xVh4ak56QI3C1VvbpIMMz5E+025Tr0bZAivU0mILSi5IrWFN0X2E2m9NgKHGkAqf
ln21osAIU7AP1iD+psdEe66sefPaGfHLCSz+0CugxLCDgMXahxQTRgno89o/ZVt/
fh9AlI/lYvJS3mV9269xii1ekd6QWJ6An7hDvYW7/TCF9w+lMCx7mU9o19yIEBJU
272rG7WX+A3vhQTbPEWoUrPN2MGfBVeVhjjneq8I4zvespLoZuIL/FZPmN6oUVpM
rk+qiQRVT5/mrcDeiT/n679c1BlC1yxw6VjMy43yqVVweu7KW58uuDx5a49fu5VK
TCegGYbd840nVCcDP53Iz6BS2Woj7SqMQF3CDUR/FKCdCbWHZCvuDQDkOfObkSXR
YpY3/4c7o+VIW+kU5CSfXBx6Nh968OPBecTUUGpkLGrhK6prSsJ9bHjL4UwJDUt5
+91J3KDr6hn7OlRxc7kYb2OPaAz48+i50UZDK4p2tNmGZ7XfC+v+T+/1g1RD+XaN
N6K17tBtDC4gymH+Ut+tyODExcD86OYjMfZZU16B0uGqTeUVlVlLxF4w8RpHMGcA
kx5AGjSjAls1bjHzNXd5wONOhWM6nG/qgVBygPyhPAI8eicpcXBG23V2bFck7na8
iTsNCrGN7f7/pExqhH35PnmRJ3i0nAKCrnoX3eFwKKCyrhABadGRfBlugM1DX4Mc
bOuxin+4xY8BA8ExBAmfxZeTECW3/LhsWdxiRxJ6QD430swIXftf8KvwGYnjAhZ3
5VMvIuu2bFIgwE7ST+W1YsvfrqpQwq/EjRGP6EeYk5WJvUIW6lYRN7N2LUODA/R/
Erz4LA9MewrqJ5k6RSKZ/2Ez0xJMqgfuiak3VZTqGei2REsPfrPCYWmnUWmXaLnS
WlLJnnavWAnph9U9+ffew5u9zXy5XkjjNNtYeJEEes5AvI3V5CYqunu4/14WqbDB
mmEXT32chYRsAsuWZ9py0fLgmZigrZlSjfdim4PpoYwDpSaMPS/dstAEaB2WO6QW
eg9ontbnz75j4BYRBOsIVOEJ4sWbRojSKcIjS/zO/qKx0K0s00N2HBlXMO5sY42E
LVZpXDDXg+3uFd258Uap688Cvn+E0t/sO4KaO1DVWrjvoIUmyR4/1PDH2h4sznDF
fdLIWwoW0/UtKpcmpTLaaZxDHfm71lLob1rhvptYgb1z/UqaTidaZfAmnCW9EVDg
ewiYq1KWMtcBzFvHYpk52lmnpuE4XaePA40WFShSvA2wNfzooS/ZsYEg4tCHbQoo
9YixnmXATe6abDFvOeboPg==
`pragma protect end_protected
