// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
MqVbsb+Xlr/jmx2CQRMBur3Ih+QgFIxDtduOrl9zPC/t4MleDiOoCjOHGtf55w5W
UIA9sSCpg6eOiWoDWvAolLXJEBsmXf59t3W6EZ5Z4l5sx5/yRlgInvFCQdESPGHK
ZVUWb9QI/MxhE8PGtoMJuZyLP8ESzzW5jXb0ZAW8r8Jdx01XSLiVZQ==
//pragma protect end_key_block
//pragma protect digest_block
EmsmrtzlIZJoG/ye/AdOihRP/o4=
//pragma protect end_digest_block
//pragma protect data_block
/WQI1HA2SNqM+uAk4xwYuNyoR/Wn0DlL1I4FYB6+iVRvddU+o8LcRUnEpli0UXhr
3LBoWJD1eJMOPHDV3Y9t6KWzu8oGI3FK84YGOQVaL9fRweGCwehFhneSaVbmM115
GMXkO549X9ufMaE8sPw9mjEzR1REAvNAa3uPVjMVqQyI6qkABKIZP5e0ioe0qb1k
E4QeyoMXySt5JHVrp+DHmwV0YJ11TfaCl4RlUeSJlgwJN8gmb+oDv+HiLauGrML0
oLGRAvzM0/VM67hfswiKYIpVCuVwee8Ox8UMACkifRcXkcEPSXHe1v6lToNV/D2C
MCkTbAWlQh6mVMX5V6hk3IROSM3zVIg8eAYTClNidIKCwnWDkdUskMl27LxMGJao
28GLzpwjLYh3FG/xWakZcWsUqPX6ZlXRwcwHzMSYF0kxijdoiSHTY4XHn8IsHEn1
sbZ2VL21Nfl4Tx9Tllc0Blg+3jCUTvXekeBUmv2Fmjid4PbMWdNJ7I2IRVEJTTDK
reotWNgm5gKq+OZxlv09xgrGr3WM2//nycrH3glN9uh1jB6d+cNwa9PLmJ8FPqxS
6OOSQPpBkgt5NCsiUbxkwBh1QNCU/Hk0abKxoNiiC6oVF94HOBBJGsUDkWOYgU5g
K09keFRk8FD98H8kNZZjbFJKCbaNXKO1qxpOxd1yTfPKxeF9ZwQULMz+BajRnFfD
54KBsD/eMbIsebfs9ds8AfC1yluIz+eS9OoapPkiYdd81VGlL9rGjdRYNEUhYtNm
8L5w+xMI7CV41nebqeGIIzNeNMtm/+K5LaIkx+kGQ/U+C/GSp4l1wSTHw/Tm8mOW
lZlN6WxyoU2Komd+/3LgW4+uO73vfU7FH83ZrYDOwonaUQuXUzZNCwTU6ZQz08GO
fs+suiJWqkCEiQuBxbSnW2qmSnfk27i6dSyoGQIMz5gcAeCaGGHb29rr+GZmaqv5
gM2ej4kXPS8eR9FQSgT+D0iYNFLYbIco3FM5QmxmScx3f0R17zAz9lJZhd6bZTVB
GfiEqPDegLNuGx4NagHNFsrPWBh7ngWhza/81EZI9dE47R2mJhQF3EzJRUqpkHEn
VXxi116aM5pqgSPcncRUrFQdYnmPyxU9XYA0emjJ255k+GVOGmNSMewD5TlX/5Jf
it0Fg1XW8TFM7cmzu8yMtbepFSK1tdrwhWVo5VcMwJdQHhsXxeZEa/cSCd/Pf/gr
Xxyswug977a5i5oD1RqcmytmLyRB1HmE/kvhPpadsvLX1gcoPGHp5RGk/WCo1vnt
Pbc+/QMhYFAYBiNVll9Gill0n7oWLGaIe2mGPjdGfS1yfIyFXqKBdmaSeNW/9qfO
eGLKrZzOtYXRXWwDfLwQLO5h5YYi2ZteRj7Sx+G4gaHOhTFnL/4Hz4KUfpXpC8KM
QYGsJl26YC5MMegZlbmFzDYy9zSnDOCLE51NgNcpT7fRx3/3gZnIHA9BePh9xkdp
KpGE+edpKdG1aQmwhuyFLsHpboQC8Z16BohMsrpE7tj9ObobeQhtSUGQU7h3TcOy
wni6dx4/sl0d2gWFhbiE6xC3M4clQz4C+gyuHLmNY5ME1hg4lFwQ9rqvc43VVj9A
xEiC+RKjd+5WyqEg3vSZFeyc5MdydQpMQawHcYdbhC1Trdi0lelNHOMRyo3r9ltM
GoOa+nizp1yiB8/e1/p8hE6lLHWe42r57n4mhYU16Z6mBj5r3/P7xd4KIMTTwF8v
KDuWoIAFYUhpJMYftEb6Yq4jS3Uy/ZsAtEPVk3ow3HQyGlZ2/pMo4PVocdKO3tHb
korouLY4CL2GHwjA1nQa9qtbYb05VFhzPLnTmnfw3XLyZid+bIsqmi6wMaX7AtKf
upxQSRHxmmqXC6+OxAunX0V8sF3qgT34PWz5sW/GJdYTvkDCEX1VFb+FoELrlwj4
S3iB2hAkMLwkT7IME0UcQV4gEB0Td9OnBmiDfhh+J19M13JyZic2PFO11QQdoD7K
4JpWHhcp+voqLdk6jtQThg5Z1dmkwXDTnT6xQRehXrac2c+B6uje6aoe+6RIwRvs
1LSAUvaoKuP5fteONqvWawbDkQkZwjlh5+Uxf6wWoXsMQOJAC1hrmZdpVOGgfKhu
ljPfaWk1J6SUcR1arbyemZTKTz5df6aTB5e2YpqzqtAVfF6SvPFLm/ouaCPGjIzQ
X1EJkMCtgghKqYgauXP7hYL5la5i1bRCAYuqDX/mOJU7MarSNLs7lwlH+MEU5+7E
rCbW6BCWIuHpsPEGPMNIixUwbh4PtoYr0oq868SJSsGC9feW0s6fkrEC9vgXsXmp
G6b8clQEyPjbftbKN4nZWBCcDzTT3QfqidlA8FvBoduEbq2TcrItlZ7tbfRPC+ON
hBf4QydXzyh3lNNfeTS3YyZZXZywQnBGaYLNg8qrJVwIaykqRW8QmTVBxS2fF1B7
bY123LrNLYWcwREKNZHhAGZD3WWHvLuHqMbTb8VJpSx1DPmGtuILFe6mV6s2jlqx
DC/z+ESJZ/cCPAljGHXa5R2OFU/DOla7E4cd7j8KCF9AKPG+kWZSq04Te/JaM/L2
1J34b+msut7bbNMLyDTO2Zrue3I5Z6yTPow/JsPYvqZhN+Xhvqg6sy8a0dBo4fBY
fQI6olu5bJukCDuCfZhexMdW5JJdMGnmlNZWKGTps6UDg+DhdWfhJ2k58L+l1lt5
wgXhpDFlJADa3Gh5kgVErofKwqO+r/UBlJi0W6lRCxtEbCZNpdYBiZrYbPzhG0s1
F2UXpyCnopPZ5wjeEFw9ULL8C8GFyVwudDX45WKUX27udFyN2/IyPYet+Q1pvzgZ
T1tDDHJQROQ/xM+QFO43TKO+LKW8TtfTZr+BYQcpZVlYr0fy1rP+Xav4t7xLaRB3
fG3na6EBDkGc9Xt6weqh/k8Ybzci1bvvvXEPqIobor+sAHyNITIDqHqs5uLe9C0C
UKEd4H+RYzRFHYuxGN7Fea02dLnP00lryABu8GhfIVlcUZrKYp/pBWhjvSoASXij
gcqWIUNgK2XzzToE+I62mg9rnaCt0GpHbuaibeGHBW03R9vjI2/p/dsRfR3C6GZV
AdEQNojh/fZDK/9xolWfSLVH2jmz27LffBuiFc10ZNQBHBhu5cdqo2PMjCbidxCb
VFbwKqRvWAkKmQPFqX/QQKO0D/n3BhfcnGD6paRfc9t8XFkpVTBrewpzz2wZLvyi
ImcwFVuoFPrfK2/tWWMHLCpYNYFC5rYh1NWRXawjEmfw/xmywO0IRyWP4/VB4Wfj
UyLXwh/kG//sAnVVABDUkj/hLq9S+snTnVDR7YT1d0XtBdyFr01iUI9lWWOYxSDK
DXfz+BhEv74/yBiKFfD5sGoFcpzLhHMMWB5aN9tGY9hkJ68+8y6tSpencXI7Vn56
K56emgIqMsF/GBQZks2SIUDouiqszRlt7Yx9QtJyPO+4CAl2m8fAJoj9ee58z/+h
f79GRFudjiJUWLTGME433GLSM3IIFJ2O8cLOZIpRNjJW7EQmNGu20hNHTygDaYee
euOKYjixbr3ybDKutS5EUUVvikIEjP7a2bV0duREtMczTrMgkFT2cyTv1RwngR6s
TxUnScUNpW8Tq2Y9BuPFK+K/ot7tyWljCwzNXYzds1OfM65JwkfSU4FBmyzg+R2N
5f1TnyRRTFadrzrNLo7QwNZO+5peAabhSRtMTKgUM7D2qEi7DDZ8mx9ST/EZmGcD
7aGCsehvhQxVxh9TvqKGupBfxjXnl2KCNdff8w7j3B9qyTpa2SjFBDPbzRPLysbA
Z1OeMFuPURF3vGTNQKxRS3SnuBv3Xr7RpmHJ+d5knoVPdQl8sEBiwtoChCxXUhhi
jhBqZcRL7RL47nFy6lpudW0TJQoyvxVQdbLS9BpUcKHKnEbahR6QUJEP6XAjKoMK
5xMN1RBy6u9zpD9WCrH/ArIjopwTlVLTbK2kbkF1HR3Hjc1+RaTknBi16pyrXfRL
B1a1w1xQ13IblY7sgz53oZ2JfrVptVJdx8ap87Wqr01YvReOETwj21zv4mfdiJgB
ha3XQvr0Q/IefR/2O2kUCAOolhPg6l2ZgXEcJu68udLCm+D93mb/fJ0dnf5ZRkld
jkVMS0W3/pFv0iE+PZx6v+V7o2yWDCpifdIyVDX3FuCJb3M8tDwQgSiM8bHEVcDM
AyAEzEuXXlNp5jB/Gk8Pfffdd9Xh+tIeaP/rHabW5k0GouTX0zt9Q5dzOVCP/OLl
tU24MSlB1g/GnJ6ZgArBFe61ZRq3UUvIk+fx3deQ+0rm1HEBjIWESWpSgPu5D1Cx
4ZQ/UX+Ru3sPokKTrZF3hMwckYbR5Mz2PUIWwcj8IJHtB2EKrcgb6SHWrZSlOVa/
A/+C086NE4At/2qtlYEH+uwJdxH72eBNPCis96MjdBlEgVyuyFJOEyUQ7BiRoLR6
N02IOjJt6jdjI75gRIND+yCr/p8FjpzX/ZQmLgJx5e/WhwvGIcPZLsPcuQBN2Zrp
3reAyXKl9Nr6MJ3Nnn4mbJWv0FmD4dRKSSWIjBCi1S1ImetsXxIV0pP+fFcwVOft
otcG4Tk6rpRxjXq9ykeGLp4xPUQtvYO1Fs3GU0mWsV+gyBe5evCzRKX0wZn0dDkS
Cnoyrx2anP9e1+tdEVjp3UEs/T7kDKp7fjQfDNHxBejKs1+YFfP6HGnTtwm+tf/Y
jiHmYzNk3jx+Vu9mnbvnETF/o/lqI73CW9iB2gpS8B74d4lZubDtgWlMC2HvrYxi
mc1zeQPcIYXgxnM8y3g/QmMcH9Pq5KcXcX8nt/0ZwOExYhZHRHLs9c0lUT9Cl+Zx
iVcYilDa1YNqPkQxtKGVTZsQOj5nAPd3YAmmW0UVbwO9Dpmk+/Og7KXaBNHGtT2H
7ninrwHIDA7kJL5fF/Qd5de5TyDugJT+6iPGPcuPfrPmyoYA7X+zRKNCAWK/PcSo
FEAggQ2PYfGkWxmwQ1eSsYeIOkK3RicRadGjoP3IG2ohZMK/QCWnnXLQgdDepEdK
vavPqwzHfEq/w/pTSDOdq/MSRw1mw7w6nUkqpGGjeKzWUOMEv4Anr0s+repFbdgh
hcJFzbf1+U8gNPqIPcLW/D/FBH4FsvIfVvSWybEo6aGgf9Iklq42HPCweHUFx7bc
yS65OjIr+rXP4hTYGzRre4owD4O7AsJyr6qw39fd3cAhzSY0XgoS+DkNt3aSifob
BHkZoWzNkPlH2hhxu0/Sndal3dJimVwtyMFBm7YYeOTjKqoTjJetljoY6jIX0nqO
oDqGOaDrB1a0pK2oQdpe01Ra6Cidvh9TU6ya/Mt5tdqXE0gCwQoUg68ydIS48WNs
HuKAhXW32LLszJDxmb1a/xZuBla27lANNs13gj38ELxZ3i1L/PjxRd8SlGf6OvJ4
ZMT0ipWRy3/+67Zo86arQY9sdqdSjPRxMkLzV1SytFVETO6RdxWAOF82o2BPPwTl
Kgs9phoQbLPCKylIz0U4oP6WMFELj4kkkj3OYNzWiG/mih4Rrs24wxT0/3jE54fM
84WvW3gqdDRzW5B1Qk+lv1p53JOJIqOdH5hzXfGT+VdsdvAA5Bt4yc2EP9qSG2PV
SQi+TqPXb5RnrF8i/wYlUof6zvgohbbqbBhJ3M3elqDa4kPzmFrS7utnkNLB/C1i
y9wWgqMQPidZypkxgPn5LOowQyYZCdWPVJ0xRk0o2xEcCP+A+YWetccXX1Ku+6Wm
QsahAMJEB9j7z5yIZyNQreL3ar9LTgyaLPUs8l0pL+oxw4S3853TTBH4jiOyF7CG
mMlqB+XyYefc8Exj5h0fdyw6RfA5KUJrBh3L02DZtD7rni51YHe9I9PdqIyJotMy
NbfP2dXjMWmwUlsrQ1t4r8TOyD3yENTdqpTbCReyQI4NM7MvDFM7vWR0nKOdiiuT
TaV31Xg9l0ZlohaELkjlKKZSHNKJPIQxUwD8/9labl3RqNRf4GcFQwexI5CCec3Q
Fm/6ydLJBHYP5XZMdMpTI1U+kado7t9y9REvSk+OLwWtuM/IkI/A5MDpI1SNm6V/
o3lQa/WFO11GRuVM3p25fa0zb0KsA90YLNb+qY0yVnj/Wam+MiV40/7Wjuq0NVt/
WTRJNgN2jJBppZUCK/RR/Mtw+6LBNvLnDfwGjVY7A0ltJcSwXyosQv1G1J/lBsCR
SiyzR5RE6Iq9N1F6SMVIqx+bmDTDjPAI4JjyZZ7PKFfEtcd5br1R4StizkO5jBXs
CLZcpYJskEsaq4V8cbV4EfntXSVil6oK1oaH8ULsJiTdPkUe5RFhu+BdhsDggJ+E
wuEJyv5QvdoNJpBKaCh16vxiyMjRchwiDwM/EfuxfiABerW9oe7pbWXhBcmue4eg
Tj3dVPxltBA0iKWwRVsF4AguO6lxKqPIpVwqhB/3+EXKbqlU8q6wo5BmZyJztC8g
SIuiMmgVFjH3v9YiW/ujzGOugUyXf6IRFrhrJLK9q9xUGkmxwRwSaXykuL+82GNi
wLL4ycAOT2eE5P9aUmta0gI7kteLthw0FhtUwFfAtw4q2HAQjre/ua1SFM/eJAd2
VugOO+wsOtSnxiIU3UkOSuEDVU4LLM6K/0Vf10Plymmg13ngmz/mVVzNJjq5HXqt
yycrWcfuZGbYuwA/veSIk5nWqqyt9biQLj89sYMGUixx0pSTQERRjI6CBctBgWO3
YYNY2nqyO+n6rcsEAoJhO2YlN9DoJAv2QRUKxst8FGTL+5BVAbPuRkymcCkL2lCD
8bFmLBN2pZjYF01AQZR3UyWsPUyDvCzHwp2AfYddG3Au6xw5rOfaRFYn4PXMjdH/
f2WbkIILhOnLwrdqN/Xf1W7WpV1WMJndnIqyDyxedVeOjVl9AyfVRk4Z6RTZPAxk
0Lr9oHtYJHNtN+LTa99jWDAoRVkuVoWUWHSyOzgxtDxvZHzvMQE3BUm0sYc5MwoB
IEZvSz23aZHl61qthOUgbm3kh+prC0pE56oVqA9a30aFYPGIhHzkHuT5J0+s0MTb
J44dWViSwi/oVRpLFVkKW4o9qsKJ+OCGMK/ikfvgbssQtYnO80wpyaZdeUCZLyno
fHNWeynsN6pj3YdDaOe+qgWTwdTzCrxDc2236Bo2lKpWTLmUXbaS1GKtPRaIqMQh
D0YrMroIhc7y7eJ1ib83sZ4CYOb6McG5QEvc/1K390BEEuj1FrFagBFDWjuC2IqL
Y6mSgLarSO3WhOqdH8l8cAvjLiMkrQGnD9wG6kStQ2qv2JR9jaGj4Ez1kKNv28VB
5C6oEpLMzxLvpgM/g7lBEE/QvIaGLwZo8pB8wjRyIggylKlN1/jG0y+SxfLmQGnp
n4NXLnmao5GqdxrTNh8+lxzGMzgEWLDoHsJJAULgUwF3xTLsA3uA9dkzAKIs7HRo
eAOF47G9GgHUY/IBDqcp095Bvoe4zcktbKKWJVha+hiVasUwfGKE3F/yCuZoek/Q
Vx3xdVO2KFR4BUawKCeP5ljhgBAMDukwiT+chl0Bx/DUMQMpUK4CPg6q6GY/0alu
u6xWRjEI3EpAPklG6x2nxCNZH5EzbOl72WnY1FhojZE6sweo71Z9FNdhJs+FAON2
ZHdmmydSJKyxrFcQxGd/s/Yb8RMs5se5VJWWS8GNfnnnrS1FrwAErhFFz47aDHDa
nFJtEUMLwB+3dlAg6+K2r8OaqfZ9kUC548RHnV/29VNl1ZiOcuoco+RAPN3ggtNR
ydBErKx4vKR7oX5d5nAIINdVwAMdgvVozJ8AeF3VRTQIUEzYnFKNsZCnbjBwD4Ut
kd+vxisBS8bo99iT19RyDnSDaqHzBQAbFiWYDRPOWBMixxySS+mGhcU+uYrFQDsG
wDb61CGvcfWLIGPuuHN/4xW8X61l9Lz/QWBZ+KjGP6/RQYLKJ1oGA07HoJ0DAgzW
6xNSLeoWPgkPZRlKAntHANgpEg77jEDab/UZCHogLAWK+WneuF8RnYORwLYRnw3U
7H2Xpa/XrNMSEXdLu8Ph5CgHHY50Ulxq9+Oct58aCVhNXA0Za4DzKmUV48rpQagZ
Ccj7Cn69alb6LgAd0sXQ/K/fNv4dh+6XTMaaqs780FTQwG1LZwvxodYA1CtTckbV
GVr9U4Pl5PAzhWE0fCN2FhfGCf8494qc8pRYtsoehiIDT0Zhs0wxmgXgIsBFuLxc
oJSAYW5Ea8rJpgYJn0J01rsYy1MIXrmgD9B1RbiiU+8mokCpbIrttGLBNhAzD5Te
3XAEPGqCZd0eAPdgB2DsSzvMccG6TnG0ivWbUlu2drKEpvyUinmBirX0dQ1zfZhX
kq+YLo2IqlZGKu0gnEHxuyeEt0xD4zg1e5LGTV3o24vr6hWk7fyAd8m3ViAnrW0y
Bj7Ikye3wxHpD8UbQ3LxcgNqNv8Ukpapdn5QZZQFrFDTCuim+8POKncD6OX0u0Ky
sxN0UkpXF9Mtr/k2ZM0gce9NcxkojtagFUHzNbKoP3Pff+UIRrbNlenwc7oxvt6X
sIlb3I7GV8Uvm60WXfuoWhqxo1/9MCkaMcaX5o7/NW2o7Sm1QUneHVexpf0gAhbd
bDD9PgHNu7r3zcmTa/R3s4pxfPlvboB+ch7mFipMeStkk1yhFy/ZmwimkCzL4Wmb
3RM02w91NOgytH0VUgOkavbXL8q3ZWWAzTnM6HntWm4eGk9i7PYixPsZnjfDU/MS
vAX1QTL17Slq+q47jGJ3hX0wrIet/Uosvla07tHzEHHS4h+Df6NJ8H29A2o1x5R7
VchG/6oMQFEsG9ohDA+h/aRow2XOpRpC5XdtxB9kU0pZ5RXPpQ2WdGT4YsyYAFSY
KKTVErFxHTX+hUcIS3OKdgLw6n0idEfXw5TEX3WsqRtPu9jq5CtBb/lhF2rvr+/3
IFm4mI5PkwsBcUQdQpZSzrO5ZkwZdlLzuJ9TdcLyCPooe7KD2SHhgx0QnI7JKhdL
G4ZzszQrQ0u5vP0w3vLOPQBxITHSKxb5xl/2imlj0IVg1RQrhe+1bC4uZD7hCvdM
hfYreTdXzdGoN0kT1GCarXUbsyf7vSwRL5vOt9tHt9RsAZHCqZb3uRjB/253Ko/9
AyDILS6BA0Zv+AHEcVvodjQ06MOiXeLNo6Lcfe5pESvkzLSZOn1scQpd7xbbck2M
aR7tY6KKiCY2355x47/bXjYk40D8ZdqTgT1KWroGtP3dV7NyKy4xVpBkdI1mFoMe
JzNyhZ6RGdYOkRB2qfNwVDb/A0cXURouofxj0VIZ5p+LLeIZ/SDTXXHpFcSRC37R
4Fe3KgKbdv7HndXTy86upMRGeDYdRE7OvTFE5OLzu4oLQGmfCu/UkJxd3g0nMZ0B
9WQFi2cpJFwGE85BBTRD7ip3z5uGmG8TxZgfAoGFLwltl8w0PeavkiHcc+sTK50L
CBPuX29LmWIym48gECw5eMFIjUw4+KYolkM05DDLNQrdqo3WDTX0kmzbWxLG+KhN
Eaeuyk9QYl31/cVYKUWMuyMUbf8gPfZHvp1+FkAJ+B70YUIh/EaOSmYSAKV60ZD+
MVci+zIFgi82FX3HaFzKEYsaxtOUquliHjkneOWe1ehYdR+11o8qAzGRt6OKYqLX
6MAbquMtbLVYpXE3Jqpxb9caPs2I+EgLcIX7HemgHfy8ZgsVW8lCCR4Tra5S8uhk
02J4BTPaiJfpAAJYoeDzVhcfqfkz3ko5380qjm9/9uxQsVezxbvJOuivX3X9u24y
G2iaPajZuTjpLw3ZNxSrNNsnwfpxwqTNyQryNfRi+CXHiX9XS2jF8Rr+FKBzr38M
O2H2UwihMZlTBvv3OvvKXnf/hbgdfj6Mbp5aFZaGKQIyV9EK31y2HS3cqqC04ZTQ
o65QG354pF3Nyd7Z6SxD580xPg5BDMJ0A4NxKUjfNNMjVdCmXF+REgoEH1Ht+l0d
apSwjWfa3uIMIuujDiyfMWgBjEZfPj4EHIBZkgCRXbKUKmDExQ2jTKQblOPVoJwb
1E1u2lA+UE/IYAOzPSn1884nGb49mx2wKeyav47Ck/P532QzVxODga3L5xYq1xHt
ZXjSjAUff48yifI3vl7uWG0HGEVqJ86pkSs786P3VdZqh9ng4L0Ong1606RqTqPo
xreBCar08auAHGRyC6vqwRGV6BFjn40EuBPg5CJKo5dMfbLdRcawYo1nUvSg9O4k
GyDLoQiLzEHeRWp6M154G+lpAhunVeJPXHuBtLL61/LJQGKr7U1pS1ZiZZpTd7c+
GOLKFyM6Kp3fEO6subv/vMjT1Km4uBk4LIEqzQ2IiLgiNNji3DRALL97cmnEBReW
veeKBc1ZeOkhrhWgNM8UtIZWSW2SjrSe2pMZXCu7HWkekRqJrex0PwnajdMp/EsR
hNH5Hvm4+2JoP52oxSecOOCrRLMfaS+xYa2y7+DigLmKCq0sXcMJw+NZbrAVnwan
/ktosi4JKlN7HRiVV59NuKsH+eRwIVjpY/YhtQZdbcotBfplO5DwaCxttafrH9+/
KEmFMH/PK2ct2o51ZIl8Ly24bMfN9eyA9CKoYhqFRudaEeHJ173pMd5mJCfno6h+
FuaOf9TaC9tWdnae77ahzeY8wQaCINhLpT3+F03Foa7txJ2ZzKvQsQEZe++QdIfH
TP7iDMGvGEskOrcu0jNQQEveHYxrC4uB2Ni1DTtWdQjeAZE53U5h7NJFSaJs4K0y
Me2mqPHkvFsdCXHz+TDT5SNfTTrIeRY9QiDP76zNKFRLf2Ej1HaDdk0h2aUfVNEE
98fjaCZhB8/yVWw2Y2YvMlOOyzSjaax1JyY9Rs/Iy0e6CUeawbTnaGCQtRouXwq8
ccwGVYc46xq8NNGaEBJQ3C9xSaxHp8SJim2YfdGystDTzEX2i9tJsTqJ/+2twIRd
gQIDXTBWw1Ua3KPtEgNWRYAdQzBR1GPrlX4Nm/a3035l0FwcobI1zdA/oMggwBxO
UkS5s3UjG6aXeyC6f/MlUWhsxzLBWmb0nAV4C/oC5SuR77snG6/t1WLyx5NtSbWf
GIxu2LuPUa8TbdqYff8yOKgPX6BL8d/Jib35k8dbVlSlmVVkhgGWa9Hv4nzHFX1d
CBFNTzAPU9J/WslGHxNlidkzhliToMslooh98AWUKG+Vmkyi04CuFevv9xGmZwHP
Q/mDo8h2l/HxRdRPsfqt0YwamxjNPa7+rPo/ZiiwSyZ6U/44EqhfX1PSPVFQ92c4
2Nt7rlalzM1XP7+JLaW3P/MnNxEt47oEoP/vPrvHlKt+UYJKw7w/OG9GsJmYskLF
sKhFxCcrkIgSdgWbMgv8eCy4Ppy0xGJGEOGlNyapf/fQvz1Yv/Jdo2hM0d3Hun65
VumOWdOmo2P/VPlg/uJ59bkbqGdRVKiEP3x4ZI7WNDLgYtmZixxytkMIxCUBQSty
5fEcJBpG8CHcSjLbvM8WI5NO9yd/bQmTE1AmxWhWRj7nx9KICA/pQuJl9nGmR+EH
WGnQOrbbxpIv52ybSemfWRQaiBGA8fMLkSZsODK0wLIjRz5zvynEYYgU3eTKefRD
FJVbqHcM30d7kaygb84W7cwPPsNWaCQ0xnVSkJ0ecBavSV7wZMt3cIIA+PFDOBKQ
hnoVXBvHPEKhiZXEwWqilyUTbtSec7oGmDmRFqK9BCzQIaSAuPNHDrwrT9TzfFiz
/M2buMFC97AsXcP1aBQ4/C3tM8jZrpu0HAM4AaSSLYYgkEgOm6poOqbHQ246BY2M
6pKyqAHfGT3DCXNx3kcZSLwsUMLWIy8zBBDOOQ5fmGOWQ7iXDD8edXudOBXGclIK
rGgdRz8pwAz7oMurmuLjXk1TCUUDTPDPVOBoDLdihKvVtrx3qdsVRvrAf7JKWnp0
i1V3V+3mJ1nhCHj0rUS1vIw4WRdDQj1f22kWXB56HFibvxODelYtI8OwjIkTWYQA
8OMA0A0sjoqSDpTQT4c45rQLLrZBzMpgbdd5BIggtKUwCu/tgjUewx+yw/N4aE5b
VzjjiD8/idDsJxtN/QZ6pbntfb6lf/obhlqj1kZpA+y03TCuby5LfOcCfu0K90Pv
GIupOA4hPMzoo8daJcvo+H9MPj1GdVmZlCvIE/wy/52JhAwdTJE6+tMZkTGc6dO6
wRI9sLslWqeYP4arj1Fo03GIDYrLdZot+qilzXL5iL/pBIbEO+r8kgVr/sFELtvN
3MT4FlsoplstX4anycXSjLg7ix4q2AcxJYUcvWsDHDZYHYNiXtBiQegjGPR+20R+
FhcuhTdmgWA+ZASnCk04IrVpR3RkbU+d/uN+2vRftsbkP6tZluKg4EarlKj3q5sW
0gh2ayhCbj1T7iqXToim6HNh2qq7RJlM7VOh7u9uf3WtaWxFvwMn3yXM/dSbG7g/
Jm4+EH5p6Y34UXQQVl8z1kZXtZdPR3Wrpd/bWDk6w2zxwUIbU3YS3r/+G8uDpOJQ
ZElo99rg0eME2B5vgY5EPmBkThbq27gPwdK4Zy/xyyNengFTkLhC4NtOJSIY+Ph8
gI9ItRMWrYhmkiMAnBSJigaXGf5KquJ72dGy+JD5UkNSv6wXIYFPjLfl3PeV0Tzu
0gnIxdmRfKjrcsqo4E5DU3XPOOsvMqwgTtgZRK3acKuZ3uNa9fad1ei7gvfN7x/s
t8MOHNuHA6ENlDmqaqUr8gjkJMpstc8zGlwT17ffrQccpOfXa6KFL21PHb67A+we
CnHobNdy3rCqxKxB38dzXUle0jOiRB9c1ol7mEK+ut2E6KtSZ+m2b6ojAPGYluXc
rkGQDFwT0/2w6a3I3hvZOVQSIV7YwNuxPgbLUOHInx3IkXjIJNLapvWicl6eaVtE
oloW6wPA23jZnOdO4Lg+ZcbXj4WzZ/CiJ1tt+O+pi6zItiFAYifO9NGrPzpSe9SQ
HZ2fouJqGkzzOXAbN800K82aqwhnJaKUZaVuyS8OC/HIqSs77Ad5kOE4ju0Q7AXi
+XoubdJ9RpHcuyEgoLhzKETt44uZm8s2vqTWjiuFAmLIx8EOXe4nIBxXPVIUaYxt
P9cF24V7EKTvtKulGFsxhbmwWsL6TJOjpJyrLMCaweylcWy3TfcaN4CTW0o1Lv16
WR/4WUPlU32+3gkNOm51PwhgZG78ZnhGj4eqmOTUluaswAzaYMifkTYPJXzQ/KDz
AqWROXoUIn+h+x2sZWQ3mrDd6lSYLRn5hmbFpS6demL4Kopvy/0ImcPylJihb2ox
PZic3y17lgCnImnQpS15eHc5t3JcyvLMrofGi3tKkQJVQqW/vZCokkXqJ+lXFLYk
382bCbuXQa/BMsmWVoYfPu0Lt3vC0bz+FzFtWbDAZjJ05i3paK+yRcU5n1w55F9t
VC3LEG7bwtMxyg9ydt3226X50y0eKhzwpBqJPdnezPSyh5h07Y2KdoGS7sDUgitc
jWaDjdBzjAK7gIHDJD1gejExm/2Ge8TQk8VvKgKxmB6s1C2gY7eNcFQjXnZyTpXx
hyHIsCF+QeNbyKtkq7+IT4wureWl771jRivWD+zE9SyWko9ElZTYjNpm65AomVMP
p3jRs+8JE9wM0Ip1GGoldXMWipyGw4KFZewFPG6HL59AdjXuolYPpODGNdIemlHQ
T0rgmCqLA4WJypwsvyYTCVy+di+zPKOjTQcnEtRc17eEKnF4eAP7GJ2yFv5OjlG9
ArSFtFKyL26CnFC+bQPFnjxorB/KCgWUYruspenxsSSI/Iyq3EDJL/hKIP56lYaS
8BiSy0rNXuOnqFNGXF0jguUqQ+08H6Qi4t5WuPUV8XzoANoBEf5AGQUQlsxTzsRN
kx72/mRDt467fALn9ISFe20koVYX5ivMz1vuoUBxWmX5h2688Bjdn3YaqnOboLTV
1eVE6oyNzmdsW3fQzcbzTJByN32M8tx23a3uKOjsF3b+qDiQnkerT7hd4+qltiUH
8rI56g7XwIR3NbxubGlpibKf5Ld9VfTdW/N8UnMwSL5FZuSWD8iE7GcxQ2gJv3PI
0g+OXZbz3N+LjJaDs/5/GmeSvfzcnInLpyITp4ioHSjkZ/eaZ5y6l1qHioOwQWUI
ne5ojz3SxNLDuliaw92oigXZRZJ04bIY8YQ2XTcfqDt3SxatDrdrC50D0c5JR09Z
7AiTTt4lPraX6R0wOqmq/DIDH0EHQJ4LD/tvuGmgPbjF4HIH6KY9N2Yv3SXSFYG/
HWbPrqxodve0jqIBL1dJBcD+BNzicf64hYp3DM8NqkJGyOnCr/fXny73GhTnn3lG
Zew5yBzpjvUE4QH1U8JUZoi9RhGGfR/wxuxn9lpl+4HbuXHsfc5MJUtN3Rgj8R66
+h2Vq+cm592gHMmOEQr7fiTmYdgZpztntAaQocy1VFAONk6FQbY5zyZDAmU2bXSH
SOPDQMi9B4OTZ60pPm8oexgLQC3qWTvLQSP+hnAv+hvOZgeDHDACZa6Ku3h7zlkZ
ItO6/l3R0zObF8S83k9QSbWAULr9pWyJrbujUaKmGjaQ3k5dtpfinVpGt2/SLPFo
xSRBcpFjalz7RgpkB5g0u6cPEZXKQt8dsKK4VospHPj8cxDgXiZAb7Me8w0fzhj5
ADIYbpjIgJ9UkF+IA7G57yw8JKPCKCvABTgDl40rHlHtmnuz4rQPIKI6522+fKRX
cQfy1jogPWHBUO1ibk4MRgPVVsjMASn9u3Gqj1eGC8zHZzK4UQ3DLizJ+/pXhr7v
sijmcK0lL/QFlJVzDThDXj7AksqghGmdXwMOC4tArsQ1R1DmFrriWHW/lulc83F1
SXZkq0FZL/WRLfmraF0sd95p+C9isJ1qlqZignC0W/Lq6AbqtZoPlK4/nISiqfQp
oLVXvShhVBk8ukb2BrUP65fFsOzNRobpMCcBNSXaf7nkl4vvJEqStXUtzRdO5+tt
trGKylBNbCctknEdkWtiUOlMkBQ3iu0Ll0m7M8sd/USoZxHrFKWcvzPAFFRjNiET
Vlxu4UWEV6P6HiuCdkgbOhZVa86UtEdQzCgXIqfjy5Sqzt3waiVukHFZGRxSywcW
tSMibPGa6/BQihDrINMjpZzQjJN25Uf70FVsjkKKjjA6bYdJUjLx6K5VQ9tOJ5G/
mCjpB0LgHH0mCQ5AwdCURHswsoLjZCX5kuRSvg89+Rh6/4Zkj8WEW9vlmstEjA3l
KSf7ye3skGku+02/EokVHwJbNsKDLK2qNh0vKxl2h3S3vpc3BfW/fKVqjtd6OTah
eXheGtm61rC2/19BsKx4tJLL6h5+CVIj93sR2nSjrYwsKBkDzUtBr1VyQ6wdHYB0
ClNGdb7pI2ggVhXfenowSJEj9kZQ2aFgwJD5S3DJtKHFT5Ct0dQIoU9PETwt/tTI
XC8pS/eIUjFvndO5Fpy2nZbW9LGZ04m1g1UQcA/7sSNVSO4TsC8T+8ai1P7jGLLA
FWBKglq4qMsrQRBgo5PlEOg8vXL394ZSfAfCLxIx9onVf2h0dosMoC99OUAHba/N
uqBSS7v2tS5UAHpHRrYCCP86dbGJWo+bQHPbvBZmWM7MaCsh4zD3h0cxw6GETcLS
2o2010Xt8b9sPB51Y4ZeIF7oxs0JaT4TtUiwIvS9NaRWjlZA/imbrUinHP2KkQrY
LKNeoFF/fb902XJhiWK1aiBvpiopMksW2cV5kSjSKivALtErYxcHlS/6FGUqRnsF
Lltuw8v4TewwROzX/uR79wb47LZUd7Sipx1ZIT/+He6JdnPyq2v3S8pnmWRI4Xif
RgVoY5k/s2YP9PXUJkVDLWVrSQOq5BN6iPph7ZOX4qzgjG+QQYqft6UNbjMew26I
UBAVjkeLfUjkHo9h0q5wU4IADQ8Tr2zNe8lClfgRsZbb86nO8jLJnQqizaBg185S
lSS4+sUhCk+1M1qSTaClzzTL6aK/xVPtZMRmHXyELZwQfC+SWpe5CJQ4ulEfEe9F
dSK0+8CdCsJ9ZGJLM8834X+PGYYLD0kXdCcFMLh7nl1vZsPJyCXPQTKxOfht7eFs
hnz8TrnaYzBqekpuF7V36RXMW6v8H0SAtVkeubgBh5Yo3cSKXDtV+MEFCaKUh1jw
c55q5a2IvibbmRZAHAXyxQra1BLmNNvV7dfKGXgTzA5H5iNJi92lmNDVNIz0++OI
+x58mpQohVst/uDyotklYEFa6DXJ1X4v8PpIdPgYJlKouSKk8dGb2DJ2I0BFkbd1
UYGGGEg4k8K6LFb4areUw7B9NtQzJyB+NVD1ZKmXpH58N294zA5Pbpfd95IQxt7v
H1S7aoYQAy7PyBmWNPQAyWxkjDYk5p+503VsuhspnVHTDdJ3fiM1tBHoD+UrDCqM
mIsEciJoHfyI9He7SOD7AcTXYwk5K7p7XHnSXO+OqAhbpbdkGqPTVxog1BQiEZui
lsfMSy/86UyHgaRYikZeftRsLXhqxo3m6T9ai5amXK2yt7steMvF76yG2XguDl+S
8OJlaFuMdBpPseY53Sq/oPSm4RRjc3I9gp4MnPZOBcd/NTmbi0ZPgrDXhBkjiFN1
C0sn/qOC3Hnot7Q3qwlDf48F/NFUhmpFDBWXn092jmAbs7sTpHkgXqUMjo1rtq7G
orRHpABEdaZqy0xSTMVNZ7FR2WVRwsVlbmHjcOmQd8doV8JwBwbEM1NZrVCX1qC9
K3GHK/ivkoK8amjVo7u81+3P3xL7a0ArN7XyXmeH4hFpAar9tbfJ5YzLqeyAqT9E
rRXcvXNxTOJ7H63kT2+W3BnkULVmGnapA9nkfHRTyWzbPaGZUVUqzY/O7zloF0Ja
O0t9k8svM/dYKdreepV7+sAMBmEIG/jC347RI3qh0wxyLVFwb4Qom55wxN7Hdpw4
0lKPCVOpVUYq3AOTs/DD8z0urLM9d7GQXh5YC73h2HKNY7Gg8Ow8vQeQFoGGTxyK
m8kRSVRUIE4fnYJeeLoQMvtQRRMz9o44pmhO7GfbYh/3MZ8XgE9PLrISv6UBxX0t
Rw9uace4OrjnMUi2vOK366mmVttR2dv1q/LA2tGBsPUxj74sHCLeIL6LtYvdb3v1
mddUNog4PCFa++JpmnrmBY1iRZ4kVbcs36ZnQrqpQtKbj/sUhLyiJiY4WkFPWmkF
NYG8qCMRVJciV+kdsg2CAuee6qwVSJ1skXp5hu86pBGhW/EUK3+XXxK/3tvObkgd
cRoyd4earQyYCxiit7ahI7eBaHK9U5qJJTNlQy0z3T2N0m1IQoJegUg4Fz+vmQ4u
lFzkR+8qqvXneRonnangnYoRG/sA9cu93/7axDVNot5bZna3L/CQ8QNrIJ+D+46Q
ZWY2OdKkFmtLw3NFr5uvpzHpkE3aeG0oHY+aVxl+1N4OxduWAspN2g3jfGDLW1Rf
GMbijUN+aM1Va9LrdyJ9ibtd2RFRi0TGio2J1RUgYsi+tuc7bp7WCJrOpv3NYTBI
7ZSq3FwXBlwe6+WxBh7nS395jfAZEXe9g+OBlF9V+FTv/+18rEg1QhyIiVLb03Uk
tuDCXURJrA1wp95rYLkvGZPeKHjol3+1RQg+VdafArktLf5gyFCOECObH5w+mYK0
XARcf6tk5rzrdSO+A0GzVdLQ10+V4o+N5Mu22/pNXrGhCMpAOPMOrrOCDTwunL+Q
m2DSmi/eD+DDy6RuvGEG7BXl+ITuEMIeC9UmSE8i7R4QYwvF9i8pErG8yk1mXliw
UuVLGj2a3wHpZ92AlKVwKptQIrLgqOA8UKyxD+IwgDuD6mOODmyM2UG1r5pJ8Q7Y
kUOSlZbU60ZaCeFiSuOXA8atz30ngdKQjSAkpqjpkygOjp1c6IZniwrDvJedXdqm
QiaQnzk87dlr1ZdwB0+HIDKf4asi1LaVxShbrzBEI3CpBum5UHpXrP/XWSqV7Dlx
qGszuioUL/1K9KMAQsDmIDhkfr0kZ0W5Le26YEc5pvsmpyOJtsIPjL1mpeUrIdJM
vn2lSwkT9J8CxOcFzfTKIc8JO+P2nix3NJuWiAcW38SI8Jbb4WDNEDCkzLo2DIRl
umYNAjikUxEcwkEulcq9a+VEi5/aUlzrcAuY51Uekgz1kqKWhm8Lr2+P0tOkGIy1
dDGMvhYVtmm8qvj6p7Z+ClVOvxMgt55pmYdpJrV8b7pgriqd/a4DkeW4DvVKS8vX
a8LCUrGEjKAafw32Pp7RnUFndpgTZ0inPBHG0fejGLFZBiqKV1CjuKBmelQODfQL
quUHAx/xcB1sRrOT1EniSzr85g2ecbpxGbRtAZirbLi+Mp9cKsteCtbisUi8QRh1
ckYBKCI+nR6qeQVVIzQf/Xcew21DJ/WaIy5i6LlYt1zlGF49czT0LhSe14+Hta2z
YiQm6uOyCqt40inIw6cW2MXhRrDPTQmeCQQmMrICig1ENSJPuHFkZxksl/Arhj1d
2dw1AAeNEx+/1guc+33mjw==
//pragma protect end_data_block
//pragma protect digest_block
ngv1nUbxfV7ieGWR8ffGtINTGcg=
//pragma protect end_digest_block
//pragma protect end_protected
