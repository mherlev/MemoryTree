// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
`pragma protect begin_protected
`pragma protect author="Altera"
`pragma protect key_keyowner="VCS"
`pragma protect key_keyname="VCS001"
`pragma protect key_method="VCS003"
`pragma protect encoding=(enctype="uuencode",bytes=200         )
`pragma protect key_block
HLAG=7 !67]A=AY>U?(SUN]$]\-V%E>%B=_)  T[!;"@>5#3FD2^</   
H[H7FAOI9/F;,EG.RRI71Q<9-8Z7:C_Q>:V$VY NYGW%, S46<A#X>@  
H)+U(ARZ7:KPV\!,ZY8]A-W0Q>"(*(XHL-OI8H.S '-:=AV2$(,HDU   
H\.9>E6C75GO#!:P\?N2<1#+I\;Z9=P-3C><ABNZ%2+GATQ)M+4(^ 0  
H%4>!V;Q)X<SD(7"PS\NV-+5:W(W4/84;=J7/DIHKBSI+3L9,KUNTE   
`pragma protect encoding=(enctype="uuencode",bytes=6720        )
`pragma protect data_method="aes128-cbc"
`pragma protect data_block
@89TUF3,HGWOGUK@\?3")/SXMC@B%K$W&J@DBB[BD-A< 
@+/B,0X8KEU+]&9@60NXM[HOC.;?[LK6K^<K^#9I+U=P 
@H+:(&[7'XP%I);U1[:HTN)@X+%_[U97QX0F%C)>UG88 
@CE?D*&&)G%Z\=;#79(CW0 .4(=B5@[NT<0'#,^RIU64 
@/O,$0*<=8BTD&5HI?FGOF X$8JZA^G+S,*GQELIJR>L 
@&?#AJIV8#?;XW$CT?_-7<3?A;'-JM^S3&-;^^MA.88< 
@]$7L>AJ./NRY0&XW[6:7>DIL/O6CSNR9=UX2G_3 TG\ 
@9XCDFYA USLS"QXMLL#]396=QHZ8T5ZS=.@,7IG]@MT 
@[[%KTJ%[P+?CWM/_;IEPJ<-J^)Z>D?OVL%.A< 64)R< 
@T-GU6OW%%-QR]NZ$)++VQ':] "'P;EQ &[NQ5S9T.E( 
@WZ3"WK6(-N6>V!<.HOJXA2)ATT9VST"'.1389,<^@QP 
@!]Q!>%I2N66YXR)8W_FK6'8[5^/[92S3YK \[Q8(=+@ 
@%OM72I2^&^Z>',UC D375G DKNE?N N]Z38P5.E:RL4 
@-3[&*<XMC!?52&H34/V=Y7)-B;_ESV<%YHL,M.UK;*P 
@U)H?E(L$>PL7(#U^8\"$61>A=&S/YW'E$?X^]YT'H:0 
@L!.T+_32?^UPO:OY@\%3I6)OUNL_/UN2=[]XH< .P;$ 
@BK9;>:1UFU]W.)=D6(G#9:^\T->F/UG(,>2.L+"E2L( 
@( )IH:_;BR!IB.%YN$AE&W@ZP+LZ<[DG92*%39NB3P8 
@=_<29]RE]>*S<0K?V 7CO:NOSYHEP+*:=PN UR\".'\ 
@)34\TLT$J::\J?DY6)YLFN'<;;SU_S5P!ZGQI05 .)  
@.^NU4$9_57W.(PP!3@[Z]2PD:*AFG]_T62FV''WX'0, 
@)ZG"WTP16]J=&3W])^+H-6LQ@@[NB(XB$6=G BR+ PX 
@XETQ//;RLFF)Q2/*5NJ  3"V=^87!/[L7"]HCIK:TLD 
@[!K-^/QH?OG J+W8^0^F[;9/UM)%!<C$,W%L:4_V!TP 
@X/2_(:)3-/6/+Z63CCW4>;H -$%CQ!EOGO&R?\-2\+4 
@K3&ZHP^*5-J$L'+O+T//8L:3C (C_I^0=$2-G3OF_]@ 
@_E@AD8H?7UWMP1'FUY_-G -47;]$F?$2%[WT@BBXK>8 
@Z8B&]\M23&/SD)H!DE"&NIR:'+I;)'IHQIR;,\XMSZ\ 
@-LHW[TDBYTZL-.MHM.$TJ6;-^,ND)]&>!#6&^K6O;AL 
@M +S<ZNQ_3S.RG>DA2=RIBQ '8!U9:/_O&7#TT8G3]$ 
@K4*7/(H'E6K,VD9:7!B(.&!#;^, Q I,A&RS .0CA&, 
@V7_GP)+VRE;$1;0>J1PNR(H .?FP:?\8XI>VNRYJU+  
@M'5P$UV@=,;IB8(\&T%QU6/!C2"IL@@.3_T6^G-M0UX 
@6A+55TQX@_V8;V[J)Z< ?H2D"4K(F?Y79%(9=OOSXBL 
@>X[HTB#9%@$$0<U!_).UB&59G.'HXL6 ->NR>*<C>$P 
@AVSKL:4H>BFEE&>\'\/^"\B>)Y=!YY:T#Q&++6'/+54 
@[H5$B'5LCM3Z6F0S:E+,93B@7?!^QGRSD2L^+.3WQP0 
@U:KFUQ_IW4%*[=YG9O3!'LBI!#);8K,1\XXV$8"L1_, 
@LCCL!G0&G_7G;>!:86E>_C TY(;\_<N6S2"W>]MY3^4 
@#&Q"DLBK_,3[3JJK306SLB%1BE<V57"BX$ *S0M,F#P 
@M 2>"?+]R\&*%CYGB(R2LTUF7W9 :?\) 0?G5X;++F< 
@N A-!DWL,+W2+%\4,7#\%< -<;WC1L!+[$<VU9 JF48 
@[A& B*!OIMDU/VGM_-4/CVXNHJF(T:3]&!UF30"Z(#X 
@Q^X @L)U(\L-@1:;AD0:"<0PA-_R\X-"B[SLFYNS<2< 
@Q0"BXK&*EE0S<W#Q:M723-AMJV0-N*7M[Z XUWSZYQH 
@P?2"<,)Q*GDV;)([U11./#;I/9@)+K>B>HNZ^O!J\X@ 
@0'?5-CI4G+3NNH8)J^ (7!$ 4@I@*Z U9TY%WI@_=*L 
@^DC-"V(]E:;SAU!"H)*4&8)$3HCQG#*N!\G,\9C4K#X 
@2!Y$A_- +1^E1&NK-:MUW3H,=2NUX"+*ZN?RKXRA,/$ 
@AO;,<O-(2Q#*?)E=%#X2TU/)IPC'*P7DJ,:PAQ5G@0< 
@$3JY;$H6(4&$'^3_!B?L]]U>#_4L=+1^@NU/CT !!:X 
@!;0$F,@H:R:PN1;F+AG1,)4XWWE2\"G#[.$",@KR-@T 
@=.7S77[X"$\NIW:N]RQ:"*_%G?P/PMV>4A3Y4&^P<7  
@RE2M# _ 0A/_>Z)>#,\=RRYBZDI@2 8.W=/N(EIL5,T 
@0';;]]C 2HCX78[^\# 5H#Q'O@- E&C!@@[F3(C96TT 
@PXR 1AUYWZN3 U* M?G8OQ%(!VG#\',%Y4$M^ZQ^MA< 
@BFF;%.=DAW3G%6 +41=6V_:>3%SD>6FIQ[<P *=R[UD 
@/K0?O-\_J7]4<]K:C>\GE6!BWDM7NC&<RKH>!M\[2"@ 
@)>4HSCYI$?!V2LM-,<X]FG%5"JG"<4L7G;X\$$^/BNP 
@-\DYNO1\(8U(RA*V'?H3[/1H?XB]ZW6/8(J>^-_E[$8 
@>8M HCT<@Q"9'\EE^30A-V\'&F&SHX:AX_:-)0T9[BP 
@[WE,!;-SQ"C&0;QYU?] E@F<=5DMHD"CI=#O$C='Z,$ 
@9.KBOV3/*V(4-114&VTA;F)VI-@^G4Y,22F5S+F-[)T 
@N_;1_7].E-!,N(P,,%D2S2TL<4]5,5-_ 4I7=\>4SJX 
@A/5I7]=IBFY$!YF>V Y)!?.PM8\;E,P@1D1X7]#NDC4 
@<6S>6G$C85B,:_;4GKWK@K2%*$CX-C52%*1Q31HY7 H 
@XTSN7I?T4I&/FKQM63_0R^6HDR^A;VLBI^I_$YUPL4, 
@/:V$BM429ITD&GJAR :>;KOS4P>X[>/P+<K;(\8.Y$\ 
@$MW7%S 4/.3J :,Z%2 S:?'+0)*86LWU;2)_S4#GH0D 
@O(\8>I%F8<FQW?9!_A)Q7@2[57RKM"#MQ(?G%^1V<4L 
@12M*OY[>&8FW^;K07E42=1IW6(S!, 1$O?"XRND4P&D 
@Z\-&PJ&Y6#@9G GTF*2[0;88T)%W2OJ4&J]Q['1J^H( 
@S%'#)F]WXL/4U]J"OZC&%+Q!FZ 7XP-E+HS =!E>I!\ 
@.C$0Q*5;7/?L"7.G)"EXB7^4G(3L>>*7N>D"\ 6 "SL 
@/YB>D<3+EI6EJIT7)_NZL^;^DDRXBV/&+:+[(L+X6C, 
@@+0B<6\*;F\,8$D'[?\"C3)$^!QP/9X[\)!00>P6B ( 
@S%<W6-S*2AI&GZ_'4/O?2;*!_D-=U&G<J1)<32Z<J]  
@FO%1.Z-6\<K80\V^@73=%>C((\+')B!3V/FH,)C7;=\ 
@]Z4D4HDY15T#+.8?%RNQ'T)=#N](K3@#ZY0,)B43[V< 
@V(;/S6-P0#JA,>:M]A1Y+/@?7O@R$\@S689*-W TE74 
@PAZ!;R,R,EUAZ)P&KO8.<VQEK\J_S@!MEQIV7G&(<UH 
@1^1WI\R1D\XO<8QP#.L,1$+I R32=A262@_B:AXEXB0 
@2U+R ,$Z$QOX!LHF<:'V3_=G(D-?S1#R\]^.26:!.O@ 
@-DXSS$2)#3?+2I.B#0AN57O4=R>"<YYN+CI+1#"<LY< 
@\AR^O?94^O-+I:6W#&>E3$(,68-#BK^D:N&&(-#^R^, 
@VU-?+=I(M#G7&?M[;7L\#ZEC.4A=5WS.KMX2A%E@QR4 
@VOV@/E8"TJP5':A!;G I"WN+R+O<&3HUQDM7+8XS#PD 
@Q B-_[?Q@Y*P[>) R,I5*!AB\(V\H[Z1(R^"BT08AP< 
@5)H*392/>VW6Z';9(:5SQ+&<8JD!AX2YP(<8-(?:2)\ 
@;CTV&O$V+[LWOUS<].HWP$!P/_]V>LZ=YSB\4GC?I:, 
@(,PH G9"L]@83D++YN^--J,^; ?EA_D\0AYC6)BC+_0 
@0?S)&+W1MU-MCMAFO\0^8\R%0_B\9(.SAPS\N]P=.I4 
@SW\X6K5 $#/W.P'FH'LO(2-U"U'=[LKKC"X0*#=5!8\ 
@0B_]N@L-X*NFKC/J*J+YT?J,^;,U_<K5M-"V(N?P_!  
@JXB#'>P)!<O&55!LDVH/%+,$;G1Q=O!0(+#98)S]ZR$ 
@7.NB3]V+D1G)B<<@AR#N3 S!6SB4)%AE]+;GLJ4E"I4 
@+AL^\82(\HHO!J^($N>>_#&$]F?(,R,KBRT\]/>:)@L 
@Y[@_=>LKD>3]F-,<?2A[TE+&C=QJ)_9OAEZ7B*FBVO8 
@(Z2S[<T$ +NXY/+?7S$+5&-Q;/*H99!=7C[91^"\F:< 
@!48B6[ '7R1<JX%C](E<,&*OI(X$=&<1SB[LRN2^VK, 
@#2+:TE,3PM6ZTJ3%!Q3M2U=F&?BXI\'X>\/+"D:4DE0 
@>X_7R;DF;,7DQ];7CX8PD\156MFG?.)^#$T6N:;03Z, 
@WJ!8SW]1^%VBX$%C-@SB'&VQ&>7J)ARJQ3: PVLW0.4 
@6WB*]8&D,S7VA2.L3ZFS>I_DGGU4H&6?ZZ0ZO1\_W,0 
@'F!#KE#@/T<-5G:HH$<C478"AK;3W3<>E80<OZSN<6, 
@.H(QL]PR1 K??KC2P_87&.$3$W$#:[1P7/#_FDS/7D4 
@"U6+6LKE.4E8! M8]$=I#F)2+"5U#^BJK=J%NT&7! P 
@&W1DO4)014VVN!?EY_GV3?J4F!?Q<K0=>35&\D4\R-0 
@K]S)EFMT_K>/SN)&!T+SN89;9,X9N(4Q<:!RHUV11*@ 
@58'$QR' >[EITVL7%FT<S14.__[]4%RA#T_@,>&7ZU< 
@X=0._/<9D":+4*;-KG;1342]2(@:O(@Q+K)7G>23@(@ 
@[6&_F@AM/L3]MZA'<3)CQN1H3 ]YR=V:X&YYB?FGL', 
@^180?TJ=>2\L:1I7Z_NXAW*!6=S#0U!E^P(;._YLL]@ 
@/C^=%DH?1,]FO(9\$P.D.&?-+?)"_3OV"2--+"/\*=0 
@R_@YQM/@0Z_<0TKGMAH4%1-!2-HR.(BFW%J@08#Z6Y@ 
@+CW4B-8;'Y-!0'H0\ZFGE2R35NKAV?QA=G3R)_@U_HH 
@0?$]E3-S=#S%8/\S(3D^.4P'([ZV\X^HI,/EH46*!S, 
@(-'A*%P.XR)(0149YALG0IZDG#'<*(91[MXZ<+1"CLP 
@&H -P1'2U#2YHXI/%]%9X?75\HO<I4YVP+7J3W+_.K0 
@L"U5[]'<EN@1C$'.[VGO@YD;1F *(7M;B&3[EB0XE$0 
@/ER.4P$FW>F6G6R>^L'^3NECQ;=MOE&KP*G@&YN)=A4 
@F1*645W;L^9JCF)U@%.%,W7KHT'ID]CEK\#1;^5S4T< 
@-%M\AGJL\5\M(_;3FD;\@4--CB%4Y:]FU%*N%68&=GL 
@HX0[^44WB;-D^5:X]S-U+/PJGE-(A'8N:9"DICP.6#0 
@XNVXEJ!LWS0K+)8DBSP3\R^"4KV8;_ZO(>0 T(J@F9, 
@DMS 58I>W->3<H8X]NS@<3S8R!7!UO:JD3D\5U_V)Q8 
@ R_J4BU<SVUV<1HC2]L$X=?^U)_DA0<@P;V!BO_A1Y( 
@)CAAH1#[HS!,6MZQ-URM7Z?KH&+%IW]MP1W.GL[.J/\ 
@X,*!<M "F-5OLDD1C*V ]2K\@?3Z'Q2Y/*"]#UG,V]X 
@C!3S6 'PWTIF 3%"L6!OS&1?4%!/PIF7[;?#F]TT()8 
@G9JP]P&;765+JWR5%XO9%VPTG$R$!#-QVSP:(?EQ*(  
@'J]J@09JG?F<?,Z>F= F^VU2HL63?F91+&OP*MC.FHT 
@#7R-=X,QN3,NA$@\(S"F+<2]6>'I*@)L+)"OK,'+7A8 
@(@*-6'R@H([#$.+?*A],Y+4M+A"P (A:8OM; /6RE8\ 
@&]VW\:]1&@?!""8R[AMQ";>>1'&7-M$Z%BIBZ.4A_8, 
@$J-A+X?(\V.%X7^,$?7+'Q@B7[)J?^Z4*YK0H'F#[#X 
@K_S5G?%/_)B_7C]\6O]M/$CU@[3>,>HELLMC 0MF:LD 
@T)<1 $QD.33?*]=R]["A^);"BL:]IU/BX">^PXGN<_P 
@#SE[..<\_W4_ I'][U.V18YX4=FKJ0_-8I%*7"$L_.4 
@(" /A/,WJ/"#/ 5\2!M'5%[J8'_;XE^XRT++IP%Q-+, 
@/^NF#LK'^&E6O,&X*6#;)4/B!U3QQ=2UODZB <67,UT 
@SX]B"N*WHS0&8&+UTB;(0[\KP;)6>B$G'/$8R'BN8>\ 
@8PV77NRX7RV1=W_Y2IBV##$C+?(M"?@^ !?5H/E(UE  
@S>G!"TR5(,X[N<5+J::3P*(V9$[U[(C$A&9E^1$-3&P 
@H>=,F C:=)X;C7Q^0E'#BYDO5^.H3!@C9)W$%H,U6SP 
@[8!"';_/]R-XD&C/V.]4 R.Y74^VSWWK"TN,A?[ ]"T 
@R9G1]C1 ?Y%=6NKPI!.V1!UP=D-XWBF %R0M[8.J)2$ 
@=P2/OZ-B5R0;)LS^"ASI.D"']3?Y4=4RIPQ=&YV#=0L 
@N(U+L?9[\ N'.4$.P&JYSBB,.1X?16K.\="XH:,\@%  
@D*GBE#QX/W@-M@?PLD>LUA(*($;5C.@XX4@5+S5'8#L 
@[M%[L4WLT+6DL8T;$.TUQH< _3JV?D(>:A!@L2(HQ[T 
@-25HB)6CV&=++=6*>%YMGQYKM#BMBF#U;(B9X9YOIG< 
@]H:LX@-<5;K!*.=;QP70D#+ORAD?Y=XUF50$MYM S-H 
@#&.6;Q: V?^@#&_-?C-@ G@FI$#!Z-AWHLA=49-8-8( 
@E:?,!I/GW64.;S:[2J+U8\/'>D#*_B)U7#@RW9;02%  
@F* P08R\70B+WABOI_D\4YW71&"6N?<(8],]W1ESQ<8 
@BT(S++ >SVJJTQ94A<&W#O(TR5:71G2PB%GM^O?YQ^\ 
@2:GDB1R@]# 5TJ<!5];?]3YAP_*O;.@LLR.)*K#]W-\ 
@92F'[%YRIO59$BTO-N99J,-_Q-D1GH$=5Z#,(6V7WP( 
@8H[%'P$6E>=8D"C-.14@%%N?*&&/'K9]'PY@EQR$S]< 
@X/0>/?*XP=-:Y=6G.U33*S2D/#6X20I62C#CU/UE<CP 
@@%:+ZTK_EQEG34[,AI :9B62>K:-M8DIA^ARE.EH/SL 
@>\A]B@B#^"3,+>UTZ+4U?P:'N(U''II*MC8':'C/&*( 
@V"L?IT?!K;PV+_?;6'&)!=4S-I[&'RLY$$U3DRU8CWX 
@83X:0[H^:_Z.)I8VK7:@GW5_'KO%<,U!*L1KW7(PIA  
@%]\JM43O'*UQ[2)%/ZMEG)ST]<WN7J .C=$4//*%>\H 
@6*&%]@*J7JW$8I7;Y/VD;]AN'=(\4\/*D':"I4?(47T 
@?.Y "/U-KY0&#%K / >X%)(P>V5S',N$QL-CP@97#-T 
@:AP5]2QPB53FU/M@<9FDO>-G[3 BV<WZDF'^Y$%(>_\ 
@]5#HFT^_I^V>H7E2['@_I]T;%D*XHA&L>K>E4&%,2;( 
@WS4]5_PR;-V6T&#$O\C?9UB4Y]]@ CH*LLP^S"D,IY4 
@(=KW2?D^*Y.I_7?TX+9@_BA%^E7G^3]0[@Z;&DC'H7< 
@ MZ<V&"<.'FO<AO$BHL^M1JM<@*=[EV5I5<N?1/P(I( 
@W_Y">=HRLC*4,H'S734[A->0N? +%DIW8(NPQ]L#_-\ 
@QPCT6@A ^B9."3E"MB7?HA?BMB9C'XLZNEO-ARSYY&0 
@>@ V%P.&0^\'^V(+1K3QB%^A)TBP7^,J2"XB8[(&08D 
@!,&-[0G@U7)Q>,22=YZ_?Q'VM)KBZ4;)B'O93?O%@,T 
@-U]Y7X6H)N@/ /NR'BGEEK+TEUS[EC;"91YTM3?0^8  
@9KZ.8C0!8!]$,E:=L>83=1!$SYI9S$'DJ^<6V"J>%\P 
@W?]4E[TR$,\#E12.;<ELH>\$SQ&5.!;RS\KE1' GXC@ 
@'AM%I6Q4ZRD%O=O8&]RINE8DUP%>X+&+W1D(^:TUE38 
@6^6[)^^=WFF@Z3%)UZ,J>S5P_Z@A=A!-T7*\RR;%FIT 
@F(1L(KCMDZXHTUDW>(5'5Y>@7B?&5[-?W?1!B<&Y</@ 
@E=*+I6Q.7YV2 T4G^8RLZQY67\-.-D'C(D*5:ZQ%['( 
@LR"#X0(%*&+@Y8XTML'4G> PY3!?G8@G=_>#@T78!<\ 
@>[ '"Q/R$DCJRMZN\0%UR.8,BA0SGG[_P3FCDO/);=( 
@>MI'.G+'C !<B],$+,[YTLD[N2FR%+J>L!K5K0G/[H0 
@#^%.5I2.N0HXA?SC#JG'1_LPM5 ]V#S1<5.F4RF5738 
@L&TT4CJ8S.J_AX4]H6:QW[*F15W2!SA[TO(F^C3_ $( 
@_70FHT!U?!,/G;?0+03'XANJ(#?B9[+B:L;/)_MF#2L 
@F)M8=<Y ,[.J?; X>;F,"!X9(\A\X""1N.KL_-^,?>8 
@R;>^K.)PZ(^.[P!#@#9'"A'1TFJ] ?\(3*1QU>9R'EL 
@00>"+.4=; B3L[@VN.?$E4Y.@8CH5<S(15%Z1\(21P8 
@$\/6<F=Y0(&D66AC+P?)<)""/B5UR0Q[-VL(0JTF$J4 
@H"?R,$L5/2HXC&\43 N/-P)D'&4K##3W3X]>V&V<FZP 
@W1SPH1&$]H5.>2@\F+')T,?\P["*I@GV*Q1ES@<$R40 
@"K_1\71G"RY27QAP3#SC9M3QN'C9OBOR%I.$S#,?68, 
@V"HUUEZ?\X9LVMN/PK4\8['B&X2IR[1QL5AC<[&J1KP 
@?D$(&R;0TCZ 8KEC$(8PWX?O@A4#)\BX8;Q_:-=#)9  
@:UL.SA6U.\L#610R"ZT1WF/?6I+.RT9WBB5O%RAIZ+L 
@:+J:V:AW:J1:62GRY61N0<2J#O5<RY+^Y84KCM2^M5P 
@+<+ZJ_K"+!.6A,.UO7;&'A0NR%F%!2'W[X'"LGW[V;@ 
@,[".1=\3E?W*''73 '&ZONQWZ>G[)'O?H@0MLM$S$YP 
@XM*+G"EQ2Q 4.;8ZYBVWNR9P&I>(BCGOJA7T*5;@LJ( 
@P#^G+EXP"'@JU=)4JPT%<#[,S#[4[8R9]."B[X^#>ID 
@$D^E?N@Q\HDWR./Z^?L/%*Q<?0P[C*Q?Y-?+1"9*B@L 
@VCS&E_PT?VBWTF7/KTK,JX-6R=J!22W>R(\CF@--4$X 
@D>+,6R4/4L2&L^O]M$O@]=]6J;#+CFD&E*6V5!P=U&  
@UEXZY&G?UXY-:U9K"C>Q5:LMWT#;A]T0*W#P@Z]AH'8 
0KZ0$X;'_1O7(,-QWPY9AQ@  
0I,#415M9T9-^VA4UCW"LB0  
`pragma protect end_protected
