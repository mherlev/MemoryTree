// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:54 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
gdrK4d4yODPRVx/BUfKvUbdqVhcXQo0bSQ/6VI+i6EOoWdEpvCx95qJf96YemYBo
y0rXAIlg9apfg5EB0PGaf0lb1i6Yq+YgmiE7iaus4kdUgvTEe8fZxpP3719yHZUd
mRUj8oqEyTJXGs/XvfCccgb/hyLHRsewrz/il+ct6nY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3232)
OaD2Y6O7AaAlkA0cGJJSyelEaDpZcRWo4P8FTUKji6vgbfU2X4ibgR82l37dcY4Z
/BWodGB8Kl5ObMxpDzBCyzqaWM/j6TAmTCFHncifj8j6jJhE/NNt6MK3I5a05gR5
Pa1EVjP3Ppt5tHRT0/Ay+J7rBUbBGrlk7+RvGsXiXACt1it6++MyL40r29vQZqhe
dLKJOMbYdrxHw/B4zTdI+mfqpMrLltG/+pKoloAUUyoeivSY0Z38F58PNJi91QY+
89aGCDoNjBVmpR02EhsCuHkxeCJn+qwWKIvTuPajR58AnIM25p+rbUGyx/IQTtv3
lifdEirRfK64iZaskuxIyhlViGO9/GyqFviLDIADGZD2122Yf3tQeoKK88TnEmDa
o/e2QIrqqn8cgLvAU+UN7KQ/ICSbz1lhU8dTnZheuAuWi1lVSXC4Qwt14czfegjK
hksrSYQ2XK1bRBjuD8zqGzDP0iOeqBvijBLzCWsWwK1pvwOuFP1R/r3Q/XHx4ld7
qfsdsCcvqZiHR0/qhhcUElhFLWiBiPvecNprvQojmdiTy3+MRwlyomjigAAUPMfw
AYx56wk28L1a13jwcbZeixdzR1eeqJu1TrQrlJWaXdBoscCGlMQSqBiWpwphp7vb
cxYYqVt8wWCuBysn3P5rjpzFPqP0OCNgcKU7LKoJLa2Ujmlw7FzsnwPUYzFWOegt
VHXAJ11BcMfv5ToJSgKKPBtH+IYcBtPLoTbqlk5nX5/1G1LFYcWzu3lyVqJgB1gN
7fSry0c8hLP4EbbDDXTcGoxGDqg2uwgLyJ5H6tJcznYZFfAeXLEHCWBecc6nzrQi
shlP2UPxXCS8RlAKLro4SslOkKH3J7keI3vAKbr1kZvoMytpK04T/5HlAT3Z/TG5
nEvQyV8a193Uxpaoi3jd2v++v5TSTXVBT0+Enaa5nyGKxeSlsBcNi4Am5aNBEM5p
meVhJv1P7gcsUiOHqtJzdGJWn5htE260Wgl59Ls5D7ohSvJzb9dPFWJQjbLpKBtW
YBilQN6i0Lhy36kLzwk46lw3UKGv8rqFg01llTxA8j2KaHO32y+QkUZ0GV+NEyGc
gBCjoOiJ3NqMEgAmnxfpdGfNMeFfDw7bAXR550lO8hfKryfV9Mf5iNO/Kaos8IoG
0kW+f2ojWQfNPtRU5jUIHSpubHUYWvw3pBBxHcTQw6mFZPCbf2g60Wtz3xvpKsUR
PR/mQ1JBfMdvbCrOZOS4ZIRZkAxXxgaYv1jQ0xTKZuEIynRZ1xK6pup4Vayp0q2i
uH28I/ja1CWyESGrUl7FivGn6q82u8qgaZHBtPzmBIanqTLmnScKKkFjXE8MkQ2j
oKbWnLJN5s6ELizflU1GEnfauabEnhXGkBPd1sErraEv5KJX8zANgeQ3cVQHTD1h
w2g1hLBhHw5Ng7VphWsyWv0EMUQn4A9nq0K2SkzyM9URjgkRspWZikoSgsArqyTz
DZTYOrzXH+NqjAPgMlJtJUKSzcHwxP883FFlKsL49rdC+r2Hn5QkvrNuiJBiFfXZ
0TpF4FwdXHPetBNv8Frhieps3Vmdhh5M6uRnpC2j1sBdKf+0x1Ae1fzYLLnQUPR0
OKwmJCsqKa6VKa01LdIZSXGh8czP61RUJLTfmiVgZYlcixqbYpw0kO5uBW9gtkcc
9ozzkB95WsVYLRl+a4F9tN3/IyoxdCostU7DhzdAtgiOQQTXNMzEiXOuTEfqPST0
LxmhJyKkl6lJzbsoIj/wEvfQCYqZo7d7OJI/UOkpiAK7uC8Gh4AYq/9B8SHvW1Vw
CgKfAEzEgCJKE65q0NARIVz4lqQTnOy2dJB9ihtp34UqD/enq43LJLChCnJFQ59A
v/6QRANk3s7aklVOXly8z1gNPNlYEoODmLnijGoh02IXWA1n0nu0aRytrJi3yWW/
sKBtsaEfwjWhZuPrvpI0iKR5r1WhmDp5HLsDOo6UwIXMwKNd0Y+UHcSYKzmu9jLC
4G7D1P/qqK1ogMmb2E3XHysNas5WsVHFQUQhfM+JCqgqeczvnEv6scwbrEz6j3pu
15B9AJ+YVMLzRD7aVzzQ+lznLIodOGPiEOtIEyZ7yB3+JxJcgRUF/UlbUTrEIMbd
bo7HDoe0lOB7yerIsNfGGtX0A3uEuDOznkydfdbGh3MiYlXQnnfCK8VsyyCDowoN
1busbKNUEfidTut8BDEX/RKKuaqbYyAr1bkUgUyuLKHcowQIIq4WwtqtMuXMbGpr
pphljhUGltZzemXmb/gth08pQ8WxUJ97GRs9qwQWrCqW9e1QMzsABkwjwEgwgz1R
TTkw85TkWToBUOtTTJsjrlPALvE8qA5alLTQGTVCpowNbVpYI/jpeb+fY+Whg1Y5
lJM41RTbExNQiuMV71aPr2G6lp/j2vP3RdD2AyVXuRFTZyrdKPYzDuNauXrquAZU
vM43M3Pjk5/bc20oEFoovfPy+S6BpyJscJu4dQYIdJEgk57bBPJCfqz3n9QhV8Cg
n1c87QImU0Qw7z9asswrPDmHLptcAGppqN1VFPuAHF6If9a+UzvxBuBcn1yIbQCT
hg+IortM6Ip5YyHE2Ptsw4d1puwxMiVbSF68TEXvY9XXwqpVv9z+QNff7yScfj1Q
IyEtIHsnyfNHmLRvsk4N0ssPd1vHFAJTK3oGjJ1aJjF2PoBk0k9L98SPylrGwcH3
QafTl4ICRSCUVOUG+YeevILp2MC0rOwn0EgfiKFd3VhidkfZGWtE2PAPlExz7uJM
7kmgnBId2bqISTw5mKvuOLD2EYGqh+0csH9VBBnk7JFJTz8wiYLnieRWjzy2g+z8
1Nz9PoeGIdNoHRqohs902cKnk5zBTZz4H1ZeZxRdXjLp/uMO9JqgyDPkrNWzuX8J
+gLfiPFDKBSLjQrqS8KSRKUT5uiabYHCfdyO/xfY4Mof3bzmWnH/pBtB1ZWAYBUt
K6SoIzAfAkXNZQTy52mDcLZ5a26G3ln779AtuMN03UnxZEacRXMVn1gnrnxj6CDw
I8P3G5HtBslVQthfWNAkW1/TuiPss9afM6jgte9rJo0VxqZ87dkucjq8xbXYBIni
RoZD3rqRfYaG/ICUSTX/h2RRob1Pnm6UKj2Z/Kx4ubAqPVF+au1Og4tre8CGkldk
/uzfbcAUvU6oHP1S5P9ylnUIGX6tSWGq+jWLdN/glkS0jr/x2Dz+iT4WxLgO2y9t
km17hAclJUZBsRmx1zkJnJurFnj8NwdC6kb2URD6JZ4JJquXqkRFVQxtXT0l4AX7
QJ/0rD+ytQF0KmddZP7YGsjrbRn3p9xRLDKepichKSBmPGy2vRVV8xJF7ihRBWvZ
XBoYdSfl9LLwvQ1SOg3FuKvW2V6zGYlEsjvH5fseaSG4/YgEyRiNvFyLgj9MTIXI
jxYWww96bbpgdRD6QT5NdR29si7Rn46Z9VcxCoKMiQ//yjQlWvaeVvfYeg6sOdIo
hrz3ZDEAuic5uqKUJohM3pLud075LCCCWaiVaX/hbNoHfZ7XJJqQ8dUakg86go2l
OX4K7am70IQuNRhFpKY1LUvucVk5UtGedD2N63GdND5r9xp2F0+GePS+aI1eqJYL
capF/fBPYKKx4rUWp7uB6+v3Pz7HlEdvkynnVNqxlbZhl5KZFaEhXxPielJ8S0BA
zcUf3vh06R1Efg6o6TaMuSaQ0FjNwO6m6FzjpZDstLYyeGubZeCgdsfnaACT1z9a
WGhCnaEKkGIlFb6bWhr0P6j5Nv2teFVg1Y/rgLIOj0TPHyTuQ0jRNkvyyq4Rs2ie
fqe/h32WPrWYqwAXA5ndkgzOdVEDJJ+IslHw5X6S4mz2gx1I4bCqz7dVU4mw+3mN
IrlGyMNFck+OQKiSXjnevWIk7t2BLJhehEtrDQwL0QPi+UyDtmiBztsJPIoupLT1
aWY6Z8UZoHx2joA25rKz96QB9C7NRyR09F5DM7rsY5vX8Eb1xFPdG2VTzk/k44jN
YnFxXR1/p/8hR/12zSIBVjwySZGK2mhB9Ug2zAVqv4NqUVnKbd9ECUc8bkuop7AD
Cz0CrxWrJoDxqZieijM6RHGKQVUhPq5n0XldlMHKNsmEeS1X62MkwdFuKXEov6OV
EjUDFU4JRGck/Fxjpj9m3hUNUMJEpmJn06kk07GsV5weLKU/bzqzxlOQFJ4bZLCj
CK8O4b9ZnhZNWS6klRlBBzgtzv1R0fG/grhN76Ral6e4BQcr0d98s5aAjCIhfeBo
hdhwhwdtKQRqkLsRXE1VN21hBh0+QF0NCpmcWzXBt5TqBQ7HLJUJ4PNx9L44xBK6
8a4kOt5SZCQCEHu5zv+ebw==
`pragma protect end_protected
