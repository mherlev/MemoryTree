// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
XLA3wdiX0l7kFk7FgKlMKyFMAdb+txH22Ovn9rVlpEsqvdPmNpWLyGQuauK/SYYpK43WBP0Mb9Gz
TIM/5KIhMw1uoYHTFdDTYM1Fr5m7fc4ej0t2qwFJsLV//CgZvuyeiNBlf2w2f/eL86iGf/9DeiGz
rV49yXlnGVzUj+Qs7raXFplsIqETV0Cdv60dxVIbrjeEnCNLx+79Xq3QGdVEFsuGGc9VsP1L81+/
oFEyxdk6yS/0Uu34dDuZZ0qp4GoDfF5maK1t4ILQWt8QFGIidHi1M+Bi1HZRaE1uZGYnIS/Ywir0
dmFcFdtI1kywtG1xZgRc9zBROfbFuq+at5wifA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
Ut2kUOHcA1/Q+IccUi+uOrb90xNprF8wPq6Xxf10p29cYyCs8tiXjYmHHCSpWE4tO6E0jEmuqM/M
slp5/3n17g6UFKPn6rNfbIOu07UN/OFF2OVTSSiZwWowhvit7407yaN77604j+D5C6MMwEYUDbC9
AXsqKc3lvWKKGWpPuFInl5FXJO4B5IdvHWEbfaLM/eNaBAPwtjvEZwnAazaoeS7aV1wbqY/3rkY1
CmfLdSSAQZ8oI19xOBZJJhr1iHNbnfN6IlTQ1EOGmMGn3YDTDXDBPt+SxH3njVdXkdywFluRmEkG
Atbl8DKr3E+bCH42I3bXrZEzN7ozJnphv6yIrEBdmhZkarMmHTGDA00oA74+mou07pwHJcyBtB2R
8lKLc2DB63y7H5JL8valDevqdXPuFqrLrGEB38Vh5BvJhLEQnJsaiBaSXtuvtD2/rYJpzSWQb96Y
a37MswQDLXylNySRw/Sc6KwgBGs7IEaRIAX2nmzZPSlP4NBATj0BddFKvouvdLWRdu2MRsR7OxEE
qFXdW6kA1L6b4yYMTTRDCaNSQpGIK9C5jn/6z/EKtj/LqgagYwJXWXjy+5W68fFOtBA8yPJApgol
jstkYV8eCyquZ7lO70r4AhJxnhwUsEW0fKr8GTb+8juWRE3GoTtEgnfMfhT/TJsd3sDeRq6h1h/R
sYpXYaVtah0X9xSFhDDaV8CAIZrw9DJ51lhn4falCKd7Tb7VJZZ9ZDegQKCbLevPWFjF3LcqpqTx
Bi7mHDVaXOTbCai14N+NGRyxEMsWpcxQ1BDW2r9T7fXTUH4DezOGExApTN+gZWpR01/VxFcbAyHW
v0gtQNdh9DfJ1NUvIZvDRDY6v3ItxOkePFtvko8n1t5Rf9OyekWVK0yDnw0mtnzBVVCjVV4PoLca
GCVb1S7v7TEZKaNOd8v6Pu1Upvi0QEH6WtARwUKku1cdwzIx+k+khA8bxwHUL7r3fd5NdddslZHv
/kRh/eQ00pou1WgAuqGpQs5AXhgcycY991x5a9SngRz+BElqT0PAisZ/3Fiei8C3lbaObW5awnZe
UQ8G04S58dWphw2xDzouvy5hFHlRZi52sTBVfC1QyMvhjHIIfqtvO5T4i/h278uw/Wr68VTD1qPk
eZVNEwZFzmWJh2o5cW1kQ74FnwiukK1YA1LikFQiBZ+6kRP+9GX9nDGbvGqDzfSNfiz5WYtQ+QGe
TfqeObT7cnp1OOEselb8WC2F2g6/EdREwT5mAILWyEJiYfihUT+0DUz4dIcZrZ7tI54TBKTF3cT9
g0TmG8LuRO40AR9bYhquEaWNn3U28SVNl5y63h2b6yU8GhtS2LRUiL9e2SXahtSWhfCAlpN4u2BG
J+UMDYJHnkb8hdctADucjDKrUKRxur93xPMlzjWkQo21FHNuJkC+by+HiyM7AY3GtTiIIQorEa44
4Ckf/GdceyboOmTteHix3+WJdDYP5GlAzF4FJFy70LNRK9WPsL5SbT5ws6M84ldXMLPSW4H+l+Ur
YQ39TlYXluwxShVDkTQoKQudcDOC8n7FHOeuM7YsyTVtswGy3fMKsMaGPTIZWWLc5u/PGKdopAni
JPpOggAM/XvqrzcAeWH0gvKb2aCfexQ75AZm08i+tCmQElqBaKoQ43hAbHf9yuT7j176Fe5qVT5+
fzGvkMKUMm2DW9bEiPAAc/YIjj6PpW409GnZJOYXPVXtoe0HYZp8jqPZMLKfxHyZQguBIEpY3ZPy
ahlE8vUg0Op1rn+5T6JwOymxQD4d+JBcfVNwkUWxOwkztt+BE9HbMnhJ34D960IX5+PcXwZpCFBk
12zXuAfivP/Wp1+fuigm+fB0dUqneIe/kSyqvUb1t8SFHWfgQ1yF+NAtArzChDGetVjke0qsiq6D
S3qTKCFIsVXqlBnHW1/zUUl/32Tg1kgqyf7KlX4jTjjZeK5tQxOSOTIJyAACma20nvVMNNxSqEiW
GdgPOnmDIoO+ePQI8MRyGD0CHgX6r07DXTnuy2QvcPQ7zuQyveLCIJhA4iC/aSBX14aRYMBdcgXr
bsCPIRpE7R69sYR6XEZucOCil9MgEiI7xcxRAO+x2bIfZ7xPOXSYym8Viha/DuT26zZZQ7c+ajod
9S+RhG8L+FdOFW3gz3Zri1h4jwuUA7yZgrg/0Cr7tNDRIKzTvHs8aEBwAzyCxBD439i7/fe4/TLP
Na7VYznBLS4uiusX0Ddw5WT+2vU/pufkcTcksyVCWeRoj0ZO8FnFUVvQdwCOnUaWM1M3/W42VY9A
Y0ZV98Iw093HX9Fb9+KOHt4Tfqgoxhm2pR8fSFKDZOypJDFtwek3H99voNSeX2hnkizfPGnILgEN
oO8+2dGRTE+SMJWjiUPGTtFiTrWexOULs208aN1yq1mkZqyyPKxLK6uqW6hGx+lXYe5BjHDaf67r
uREZfz+ZsqUBM3kIvruXkcUDKMQ3nLXV3zjFnQNT9PWwi5aiJWv59Lz/hnqSLab71gfTfkIpz0vJ
/Yx6VzQqYjTD2MOxilvV7Mn6PbK1ZAX3ytm82IEDqq7brkXIWO2NBakBtuUQ+KV9pVpJakMBCP7N
u5n5E98ShdIjChxzKUwlvEi1WujSEwzYRQ3+R1XB0ChjhgENcT4htO2hKmDKsGNQhrAyANh5XEup
tTaTD+Tp5HbvCkbf1pcZ6xoX/w/CqHGYitqb2fiKWazV6HXewYdt2C4zNHKIB2pgAfF07rrJ4/GZ
RN7w+FCh3OWFKblIm0pj/3igIxhkHL5FT787T6UDPcKV6UoqvcjIon5TTr+PzihgxFpkrD7ofk84
fMa+EziZ1j3GmE8R0dHujj6sJ9TP2jUHoqAwe+ZGsO2CDBl3WMEw20iACJWS0136CeVKZhE1/1i0
OD2JuJVK6RdeK9yESrdsgbMeKuEViKR4tmjJt6G2oF/3Dc0If5fMx41CVKbQQZCB1apcCSsyBQn8
WkRp6VCPQdjqKtpEEEkmQb9pM6Eln3WSfVEPTYUxVXal6uU1rAJeYTS56dVOT909ni+SYjXaYCQG
qbJA3ZfaKe5JsayGDictNKiZ/BVQT/BezwhFnqh9mQdm6RiUSGYFwWoQb/pNErv6bcYtzEd7Voe3
nHl0PjJXEl7DDSCo0nw1Fm5oTC+ICAANcotpcoQ1vyxjupWhEdS+XCXuoED+NrfGYGjmiCFB/O/B
qrvbneLRBUo7MFhqr0QMieCzG0JHpgjbTTgLVYdmnq5flpn+ePlqTCf87I3qOK8O/6ryn+5/IKlT
B732Ll0u/k0EIWDUO6j53+qDHNqImNEPRsyB+lFmvy1tNUwLQr6IC4tTbDcCaj2B35bxUSVOotY3
juXOzfl4n5x3/FFcQkbxPmUakgdy5t3XwCiy0MH/vOOBfXo1cFfE2DnfZSU4L9FH2ZA53HazifjE
py2oSHoUazOXvd5ungF4b3071FCzUznahSZKWojOMog5r8OKFTTCFuXlyxPopiydFA83ji9OL2Lf
PIkofewOW6OSLBhnn8WY1vo81kNI7Gr906WnfjcfiLciSt9A1B9C//ZySuDarwbHssdl0EHsOSyi
uUmO2UkZ3G4YTCkG28htHo128nk2B0E7btZ5cFbSYf6Yx4VZ7svzzx6H4yqxxQoeC3P6CaWCAx0Q
JpR4gB7dHQ0CE867x8arZrJuN1SS5ce8qyPssbv+wcioLiZDuFl+QarAW7CI7XFAMUKyjc3On5Du
qFI5hLQ2ibRTGdjgH0LCybTI4L8WWCzf9JCsZrJ9zqFuiTFqN7W6BHKcY3GKNkCg0gziq6hAhBOt
q+NB8bJiqp89gKa1GxNPDG++GXjN913TvqPAG1fYv+MKoXFxR/PDDF7F+JM2b3vhRvUpO1hZsfaP
WJU7jPE77KN3ysL+wyjVrsy/q6vEUBDPudNm2J5A/z+a7Kq636/twZxgYAgJ1SqxLWRScoG/htyU
9eWrfIdhufBj+lMUPw1y9pubk/sKM71Iqi4KBPFJCikyK4gIaATnAx+dCh+ott9fN4HRzYh9TLJG
NLfEaeOrnYwwEnQY2epvUkiN2QDZbBu0PCjpvhICp0mpFLaBKt2k7votphl13dxyYETw4l2T+DzT
MwWTaKpAw0j59P5/hLd16bD0W6NJ5iDcxsn/Ij8xmxmyle7jxcHdbXyHyQhKpWUwC2NoOFaXboux
JgtGGn5IOj6+XtopkrBlcYbqBjknTgChJqlA0MPUd42/p8l82jr7KrpjlJxSkwEH4du8k4vxdkZ1
GCkbcqowxdmK1beLqQrayBlIaVZOc1iEqWp4pahJoG2djhE8v5UvP84A8X6tj35mTk6AAM0FOO5z
BHc5/MEyMY5KU+x36ZjvqVSMBoEEjPadbgEZxKsPhhI4X4zU/iQLvBHOCvLaQ2f9hB/zOD/78GEX
3VfSTLW+4p4ZJo8Q8a0JlJxYxgs/28sg34QusHY4VHzYunmZYjqE5x+vk458PS5bFd3/czMpewOH
iRqB5tGD6t/xSJIEqKj5OJHh0oziWP/Bcjv+/wHBLlXXNI45+Az0GRTIQfyErk2M24Hft1mpQiUs
E5h1C3gBaQ4e9siNs4dd3EkmYrb+SfvCv0HlpUNB84dxBaUh1Gu0X/omjtQ6gxCRtRzI3nVcOnk9
lrgC53U1lpqUrUmnxIQefLhxjZK0+XHe4im5S/6kF1rxaNe4/PCVjE6iOlCM6c109/MOMmF2FDTj
mqQK9Pc3kwBN0tzGqH0j7nsUgOkj61gkzasNG+/KMnKk8jMUMqFPu6GaMsJTDX+0cWVDhPArs477
/ftEazQYLJDWo5ZMkelIj1SBiwD5Sllb4uicCsT6ZxBl8RhY9pN8b0NZLFkVwtnFC4xH7Od1wRi8
4+bZ7a2OEw15FZpJ+rTdZtIW0I+IlR7KpSUvNGoep1dL/xZZ3io/ootybO9EpCwVzRWzLJvoioBc
v51e2mULDtcUeF25AkoMLmQuZCK1VYeYecjY/I6bCRSyYgLpyB3T+EC9ArbUtNSFQJ2bDUUorKsc
WmNB8ye4LzpZnf2xXrL1wX6+bi+izIg1MF8ZaDr2rWgFGu9CmwQpcGbBXzEsvtmawnAtIh7C7Obg
6HfCOtq4ID2XE2yiNHeucde0zeWffcpbTFZ8VdSHRar6ZjYHUlaBbdX7AnoPYDRz/Ut1r4yt0Gvm
ekoZ8T3w6rwaTSmWTiSg+44Rc9aXtjKHyP3HQ/YScgTUwJslDb8BBsrfaETzAF5Otkmmo13CwJqS
nMulPBK3rv6+7Cpz15U0o+7LVEIkbhkiah/ppoiBv5us2sDEx78zPacO/sXDA3NcaC2uWHubD6Wn
pzQV+0rq/dVM9jqcUPyHYlcvzG+9l24H8q6SrtsP1adAQR+aiY621zYgLIdTCURZqDXeTGK21mvx
nZAnLipOJ90ss+xY7XmHMVkPp/F7LB22z16QSeSCsB+fi6WouL+JYPaFL+5tL8doPLyNwOX8yYGJ
tvblWWGUQ9MKj21GTP0fNqjvucNObtrKXjeKVHiBswPaFeMdeXUPkvTdT0+/fOMmRe/OnWedJ8bm
orkPu8kRGQpgD1nQX7W94NZee1B0PjXG+SjCGT3hT3gTZbk5O4ozD0I3X4dghF5iTq8CD5MPlgfQ
AFPS7iucw8tT5YP38oh26XXvYkvVs/Hdu0i2usG+OkuQRJjCbuAhlMQFZTbKEDFSv/wW8m+sHIro
7i8hbF9OD0SsA4U54ElFeBUysHXuCqrY+GPLk0VQkwDCHAx4wUN8QRmoqmbTxidddEa9IIIy4TXM
8UHjRZF/fAtRymsoSL5BsKImJikEgcqDEIQo4DLZHuJopKK03m7IRFyjAXlqTXdpEl1VSMGKg7f5
wRWEh1DsV8ixvtsvR0XWDicb9FVbbZNBTDbIgNc5WMvEG8Lbp02dbpN1wI91wsX60QENAnIy50No
EAgHGePTITPjkGwMwrhYW0BGeHJQGO2MNbgG0Gh/hpirQG/uFUhboLxZpZLJij9cnYPK4In/g8fY
C1pAGlzKSKGIT6u1iPYa4J4RmyGNdZZ49NovzdjKw05wQktX2obFrZSimuY3NXvyODFfFeAZ4MzF
CaFNzxF8iBxHpbhz+KYmozL2lZ9t+LfLg7inndSBaSDR/G9ccy31rA3j/BQ6Sohy5OpebNsKWB5v
V7Gjc+yeQx03bF+HwyxOA64EC4h7i4wbIHJqoYqzowIytC7crv58XA+RMk+yxMyAtAvfia5Zrr9r
flKJaZYMLQJyEXZh57YAQfDVmWgDLPCebjIyARbLNekpueNV+FmSwp59CPpj/6FI+jDEO+WBQlk/
/9IREa0PfaQ+Inq1qvR63vOtoQMSWyDfpaxXw0xAZokUfa5fjenoHqPkOq1gWOIiWSApLoMsLvpo
lPaRrE4DgXJl1OX1lIpBtC1o5Ms3RT7oJrxbInAcBVwGLtz25ayFZo+w18qW+Rq+VtY1hpB4NRwm
9joUDAvceu3q+f6XqvXM5ZLTNJsn6DjR5aLvajL83gcFdHc2Y4JpnH8j81MCxfNtdHYHWiWZQj3o
UeDdUVYxxY9nikbFAa/+1AWmzHoGIhGR0cfbQghZk2yHqXiEJa35+1vMJlE7vv4mUJ59PvLGS5Pa
i4fOueedkfu0ggGcxKbIj3NmoGI4hbfhalVyvGG9WZodxhPx4tiS17GIv25T8+sqMwX6g2Te0FyR
Z1YQ37MWJ8rs2l0aZwEyxvTpFvRh9FPJuPIWfT0/L3ugDXupUO7LeEDp7LCHV94+5/KcI47Mlspt
USDepzbiGMgBZH0UXqOWaqIrH/3xPpfEwdp2J9AXIKvDD9uHZyOxY/1p9tOr+lzFI/kg5n1kittB
fwzEZ2adazyRVrNwevnJB4aaiGc6kQzxip/DXhi4crTNzf1y2cpYWllWcg/DRn43RSbwEOQfocKQ
5bk6H2tm56p8BiZs/UgZaLlZt4j4uM54U/6pn75eitVerBOr+LsCXlkfZEt0SUzT1K/1eVPZrEj4
OQfyj87LQV7q9EkFuNN1LHIONKTlj7BQa2YBrCS1tEbpLg90WRpfXUJ9QPb8m5+N4uTHS6UVJqUx
Sl8xkdZgpuGg3N1Zo1XGOukFWCyNLqvocy2vzfebHmxFdjjYbRWDgRrrVU/fT0Outh8PmjvobFaN
xLjjXZUMwrwXRnYDxej2cb/wKLyo6oauXo7scOPTeRHlGrHmIZDU4Q50+kE1VVwjxcNMYdOFfPDd
rE1gcx6ERODr5hg0fWE7CPee7bvbie3mtEqP5fOFuEMx6mU8et3o/hDUyIFzjYlbWgXq4Ubg04sp
uPTSiWowpSt+a75Fw7xyqas8OfTbJGvZbdREiL6lZQReLIuSVTNmzkp8XGIdE8sZHmZVOtjSAd4r
a1IY2ZdithhxNdCxnYePbZRsiSt9GjjYM44AI1XaK5DkCvhuzuUSmv5sf8DusJIgR4gDClePA40q
IxOB906jZSWJPx9+OJ/d0TW8C3Id3Vtpjw8UsAAcqVuz9xFyokDxZviU7f0rOJLsxwCfltPZUsF0
sIpcxV1oOdlmFi1A8vSt2fQicpAmSYX7Ppj3V6vF+1CQ3PkhLQdLW1xLvTCPbHTkPwTf4al4qKjN
ABPVap8cMFR7C06x1MEaxaETFdLHfD3m+aza0kO6R2qGLKnDJi/irccTQV1d8Ox9odVa949EZMUW
KvsgdG97MHWVnAoexLX+vQHvsuzNzsb8/AKTw06McmEZs6sICeBVeJgRxgBjh7EaHI1RXcwmjXTY
Ujp03KhMupIuQzmWuX/5yPKRYE9CEX53WRLhhX2zyJHhYGPvoXnUf/zGosyUolINZuHZbg5sq1JH
sx84zlBzvFVmzZuNAsx2HngiBgazOfEm+jpqhFhzmpc7ieIS7XRM11Hg01NVuibinwd0o96J4U0H
sIKYMMyfwwpLT4HmpcJebGOjV6nCOMZzoWSdpAtiPLtp4dfdXodXokZqovD1cRl9IbV+J3VwACoD
1a7KV35DFA3TbRibzYTwNY7BpcwopeMHMqgNODDw1CfdmlONesPDIj+Tm6353myyz9kG2mKzUTVB
BAv1Kjs/1qfd6wFKd8kTTglMDBh31jbVKj8boVYNrr43V5jSpHFPaOhm3TVCowMesuvRzQNYVL02
JeCD1H+Z+j79Ly8aF6BxxF+7uF60b7ladUPIfrNhnRGVJmOCdbtUFceBMoxd/la63qjWWeTeNTkB
9dYKsihVH8dSNuAoVzAm7fKKLVbEa2KooL3z89jL8BLavajZXBbUFdbbXOQdv/Ty9NYH8WqjT0NH
6ygcdw7Z0V/WCW26Vv+Y0/LBGU7HDvokLG8EQ7yHv3ujBSqd/Gkn/K0egTDU4X/BoVzn+F9yT3fU
gA9PkR5hFBBt3IR1PT4yCimlDi6ZeJMvFHp4yXCRWQYxWG5kxRzr3RolkpDfdRITchO5v/4gvXAf
VVzYoxBMm2THS4+Nw0VUo6MSpYBHyqbPVXxeVsw6byf+R9x6LnVYNpTEH+p2yUHGbj1jc6z2KSsU
jJf9evjTxLnLVVsJgPQ8/RqQ9/fOAGwwewwXWYi3yIP/lsIQyWwbw67Un9orAs01cxURwrJJNzIf
+j2fh/Rw/LBiM61jZhWT4z0wcZHjkMCMYwPCRKcPn9pil4Rwnp5Lw+hRiYM9QPholsWEwM0YPYhG
FCF4N59GAS0tORMmI49vsOOSpJ1pUlE9shCcJVW8cuxB3VeOTHWUIBEj5Wlyj0UhwaQpcRH2KKdM
eUV24+if36Cy6fjmev1NICisl/Z0KBZQhIpNFvDVT+21Ur0DAQdSFuZPxUZja9u0sd7BHnQI1vOE
PEejGp5PRYqyZ6ScBuXlBBGU673czIVh/zcJhEti3OQnQXxS57PTYYM9GX1WT/4PosmQlL+EnCmw
g97fRBwjlhfyJfah7fK+TtsX0nEDMVNuw3B2uBakbPAU7SLunf1X3w/Sawi54V4XvHFEcHjuncnq
f6UpFynYJuIrq0CrU0sKYHNEItATDyQ52rp2L584fNwBiFzrOpDoyHxqEUY/qkXckukdVO5fRls9
oes5upDkneCqucKiuO5mZ7Dxqiqp2SAFKnpiQ/FU1Cd4M5kmXRoKKYqWAgs0VxwLZ73ZtwjPWT6/
RT0L6PfBicmySu0eZbeBnI2mv91Og2yGYf3jspZNWfmprnGVNfnR3Hy2jeNeEUe3+6a48+H2XRJh
oq1sFhHAR22NFgEwxZ3L1qHvnp81/LvZwVL0CvsfMhKdcQUJwC4ULZ2cmaDTvCZtHReQTWzz2I9i
JvIcFyDnDHvSnNedLZ8egpF5qwzaCRGoXWTmCwyULEEQ6EuVjV/97CV6ykhL51zKsc7GG9CqYoyG
olctPzlTFv64Vo/uX/TrIfV+40URNXGJ4hTPAmL2zZA0UBprDqYN3YBbDK+G+1uvwpxkgLcHIKWG
HHZ6RMRmAfwjLAZD48VkF8/dwaXq0EjsdYa+jow/qPfXEb+HrgFr3yuuLlhd2GGd0nIeBTQnOa3y
txN8tns+QrjsWkGILLZ5pNqWhJvyfydxmzlsY+Qy40wWRSFLVp9QEWxdWNYSEoiEAwXbYdIEcoKs
ZEtOPLbAn0QgzBuQDvdM6agJVxTKiJGa71tVN/4Gi4cLXzDo7FR34QvBa6BT8CvtFYIEKRk4nlBN
CJMClcZRZVIvdWdoSYRLy5gAhSS+Gfol8Nl+nnyjKv6RfolIQygjS0uTn/YjszJ2gzu1es2REMoI
wZ+LO5RFJHLzY9lD25KvH00te5nDZ01Bm6UgLv2SxVSdaPrFH9H2EGl4zPYRJuv5n66InvHQiWh4
QiFjEaT52Ljvr21V8gdVxJPmZheCVXaaL/nBABa/LPGPC0DafzMfPFgNo41X3kvTU15aLcNQGfqN
3+De2dYs7JLXqy4AnmJlHynmFGGWZBzkHCATOzGxkMq4X1HteRvpRWuCJcHCHCL1E5anqEi8mxRz
zgWRpWTe+HFh7A9PNvLcCNIu7qGPEUuwljlUQCT+96QF2ZTzA7MvOpNaCqtX3TqsAhpyWWq30mP+
y8GC6d9GzfHJoG25RLBGVaA+Udrwh1sTq+3ae7HZsf6KvHcetfR69fxPDoEGbL63IHM5JJJYarMG
RxsNYmrclYn6IdLH/T6XrEFs0HQgbzU3reIZLvml2+XxxwmN/1eIf92xnO9h3O3QhiRFQ3wWAUtC
80L5SVAXrHwC5y/1Jlg7nV5S6YcWh+Dqls0ymzPqoPl3Yu3nrjmhQ5PNqFwuHKGHfjbUAo1WsD+g
QXX4FpFM8cyf4Z8e2lAmHdqmkji8UH5cVqDciUauF+yFciyKY4/lie8TxQ9WyRjNHu49WoxhJEdS
TRvBXk3rl9fJkUZK6wbbb2xHR7npBySjnaIZQL4ZHmJgecCwVPQGeGbBPKRDAfIIu53s26j1CatY
C8DsQS+D0RtexWgG92kHvKmHz51zgoz+K4VkTryjDyoFoAeXbpOswEb7fnEsdCznASh92T476WtJ
n7FqRLf82y6we0vYBHI80NWpqOJsZYkRNpMXKKQ/eCDVQMBd3oGyNn50oPxLN+TDoktVnl6qGK4L
0wLaAhOOofE9VKFlSxwM7YS94qok6H07SboJX8aeAmR0pING1irKACuBQu1ZUdLYAjdaY59pxay9
+giN7MM1TXTAC1rBjETWEQj58FOu6NIldbSYZhX557Fg7awL7bZHVC5UUHq9MDGY4aiKLTRTMUbE
UlBHxlg7uzekVWJZ7riy9Jc9fNCPiqYh1eq0BrwGHcWi1rPr8+tfNCncNslxsVd2dJMWdlRSTWce
t5EQrQQabLFu6d5X2Geo8qsaAXeZ9QOra9LKD+cBlVn0QzShrMXoCKYAGDE/Pj6qUseTEHt+V/29
RZGA6jWHPe+5M0XxdIc5+S9dA15+VIkNMn5Y0XYTkRGdYnkHrn+Zn8pAnDZqALtmF4vypboyMjNx
caW0WOLWDSpOUAxgG3Jchn7PaatLAK0INhHS6G33VvXQIJ43gr+kVKW2XN9UJlSZJmyiB8lCveOj
B8FjigFdbYTE0U89zSWZxNnFHOJaBoG2mh8KKOytYrgTJk7Hn8PXK8VCdcslXHuiacCLCR2k/VDl
L4rMkt7fxiYTJNaD2u6O8YlE12vI7OgDx57n2qrf6r0WQkwfq5hdQu3kakZGKOyg7XpkxdYDeszk
RiuG1g8czrduhJUudDYLrUSVWsoC2KDV6DXSCIxx8dfnoAq4tkaURHWPLXHy3jj49SRUpCF7jjSm
crFAVZLTu/LcZlaqCoXtA+eSnLNgrnYzpH8C+HP6EOHLEUQI448F4uR/cxS63iC2Bz6dKOinBw00
Uq24ZZwIoNSzy0Azkwl2m2Fpp9zjPrai2qg3r1RhdFgL9TSr1YVh3kZIjYSpezsjQB0X4H/Af1lQ
n2j7ElSpV4l9WKXreQng0+9pTPYgQ8sknwKgDvFjYxjGfCckcOzBgSXYjEPsE45wC7RzcAwEbDFp
DYPzTPCxNLwjvxg8RY2MyGK4jQ8oGbOs2arhy6LwnP/V2WkvHLPqvQIKhIDWkCXdlvZPDBJLv9hE
k+qV71lmMQeXSMwWZgn5AK31fKzUKM0XZ1DE0PW2oBqKBu84C6b46A+kSEHvEpEo6qgsYRjBO8V3
eZFDcYY+bKntGj+YR4YEz9jLda1cef6AXl2hk6MuYcoiofOT5tuEewFO1NdabXxuGnNpspR4bABu
JTezWucd5aA2/4XKIErZMpxbqADE27BmSICBdIYHks5bbGZha1rEvbK4BAvK29b36w3Lpm8CZGiI
noYRujv34lx4FeptXgt1bMNPetJhU6tZYX0oWtabOf8dsAg91OgpCts5h6kERopcCU9kC7R8fKdn
BIrq97QKYbitCLJ6PSLQ5uuTjpIlIfw4CqNHPWv+9KIIF0UcszddRQVRpymnyPnwDzhdn2MQi6MY
ew7qPmeXW63fDlu5mUP0/8QM2O5VquOUdiO4+6UWSF4HMY6UGVAVnnAx1Pya1f4CJGTReB2pmmIs
rdh0lyf5pD15dIjx6OSQEvsPGxIFigyY6YJPJA6LbB3+gxSDFSzVw/vf72PhugZFbp22q95bCwNk
mXYa7v4p4NUwnGk6mx4+nbdlk2OoqsWYNDmc9lOr6+TlpQ3BQJcJYOppa8sCWFUB2tUFa5KWkh2P
9p71kVUceY3Dwb+nKofdX6Q9+WQBjFgd9KFAhrOvApC67H8o1beGVR2aIaxXpkY4Mugiy0b3pbVW
9rFIOobe34FCcLQLPQrf3NLNh49xuox2V0ZUDJxXe5ajXJw25cVhgodxNR3XCz9co2pAOMMYF3zI
h+x3vEm5+HfJYUpQRVihpuUYVK4NRoPp2hM4E7NW+LS8TFv4iAbPUedaLy16V8oLlY+ieafR3PXp
/j4iBf8fgnY0mMdMxSY7FlNf5JHLg1/xS7c5VgZ/SNpl09OqA0LlrM7lCSYnAZ2uWcRNPJgLOArE
B9rDgzuz5m6xhmuAdS7cmWdAtklsVwY4AVqTLGsP8XtfOq/4EKE1shCZC7Ix/SFzmOn8KC9UT6Qp
JtvuJZEEQUyFZMaFzbXW4vJC9RblhdDi/8iSL65r3ijcQwVLMsUUZ0+XavJWq8mf9wtb1bGKWpZW
KIUpTrnOZGfEoVhOUE48/TsfacrCCGFAi9UUGmxmowO1rKI8kt/y4Nkfl3kYjuLzQUJdBy2fXr8M
NPQ0Qn6cqOj4am7eMlqU7secT3S7f0oCHdBURaGLZvNIOfBcWdTYg+6RK+Sp8ekF6d4bekM7pGex
m+WrC5IX8uLP9CeTYIUw9Ajn4OBw6PPWHOnYcU70g5uuh57CtGQaCPPdRIkxq+j5VJ5cEJAKWQuz
8dDTFkn30tGYwzq1D1aA3EJO5q1IpqjZ4FRo0FYI6uXWrxfeRuFiYuU3xpstyaDNKHWlAa5twG/r
g1mNRsYyJdyraSYrcY3G2MKgyRuiE7j+wOODp2mwnT8D9vummyrGA+Bj42uptRn1mQL6FNoKgyGG
2F+ppN5kZkMGin6hqNsVlF+PSbTItc29wrMco1hU4vSOIOZXzlhc0eefOLquowk5FSTcdxivv+fm
aSQbaCvrdIZdfWbKXrX2fNgTBLYXDsDMBYmz82LKj1RkARVfLM4WoOBcMCK69QAl8pRTZ80KEWgh
hpLgRPBJovf7X8wM+NYAm836bogQIEUL3iO32U/kgKZBTyTzBMoCVjRmu/peUvYr8PVyuW+eHAvk
d9GQ3t9gRYJVTwhhvMO6j044rTY4eiBoANNCyW8ehzu2o2bFMKS/dSETriV7Kxd/YXaxu8q+FwIc
qRPy/hy50gdJRqgEc2A7msw5As2/qmHxVTqy5kKtg8LUBQrCu3vwiCYczcyoso6ga8YFpPMVcpYs
em3V1cgGKG/vv7F39rty8Oi2trfqtHTg15ruL9qENQn4oY/FINF68WCmKlpr4ToaVmP2Cet2Ulpi
Iv4y8n1i+lohG3fPjU8IShW8Sj/ijNDzihs3CKpNspBDZjxpdMgy0qKcwdt1el/Z9BNrw9224Fce
77x1yft33hrLl6VrQzeBTK14/TpQLyOAvOquikDvgaLtfvHW69QT6OJfDvDVsh6fb+vYaYGNvaTl
Ys+uebDDmijO3ZXwBekOrVsvSTo81I2vnyFaX/W5CVREjm9A7g3oz43HJZRcZjutZxzQJs0JtXCN
PwaB230harnCTok9tDbCYyj/9r67JJ0Sz7y/lipcRb4iBtIlpboA9pAkHWSAIqDzX/TjV3LilYbL
4yVaklRFwWdOpqO5xhvSv09zx4e+gxJT/J2/95C5IC6Ycsp+Gi/1t4ai/6wWznjzNNZJ58V9Uy18
b9zaQ21r3JIwm167Edxkkd7m9hrTJkO8cLUzlrT6S6Y9a2Q9xWYNB2BjHqfk32R7HPFRDgoupACU
UUcxeNfhvQhHiuVvXN74v8hWuBBlkaXdJD7c8BV4wtiDdAPc3fJXnVh9PBxzTL1jifDwfntoY+br
TI+Sr1gQzqpLOFh1bTvU2xTEQGqJNmfmmXHu17DOuZ6qnWkduQV6yWXXJhnyg6DX/Oef1ygO3PJ3
riL3+F73RgDQMilV1IAsOhYb2ixJqZDGAdTALPaKApJ4Tysl5y0PW3wlc102etKlcjvaM9iG4rK+
etyUiBKyv7104j3q397QX9B1OnpW/+islSr5a5TfkluRHsOaSjrsWbeVaYwGFWTUKOsw9MKWT2NL
uJM+irc6c/Og25unUBewSdtyt0W/jzgmjcL0NJVODaAKEjF/habV8fVH/mBbgf5N4+vouGYBSj7a
p3dNSDlMdiHv9BfNlEOeQtOByeDlS8r5kFbIR14GXh7vrMxiAzRy00yzR7PC8jn1y/y2kA4PiYAZ
+LJNN+CFFM03kr7cXjyEgJkFtfO7Ea0CZA02jn5FZrLlpmS4KJEmW+4VYxGVL/CXONtzp8XXEXU6
sZyWN4x0SHJ7GewyyC7fWFAn/advYZNw95IXGsBFcSP6PTQF+OrucldS3DbCkXyKALcvW4lKSeGk
m8U9B+1hqj0ifJVoP/nIsTTzrfkyTURwDWLOoIjcWrjvxzjstgo5R8jWvLiQdHMc6jLgj6C+nSP9
hRlSa/8xa3BqkM+LltsqHs97FV6tvokVU09Ch0s/2fgPjss/Jo7bV/tKfuc58ImIqzgJ7uftqBam
UkVw6Yuhs/BCpDM/f7wQNTD6rFaLZTXtMWceUZfpORLyWvuLNTkp8WuollKTwKLLRjlM3Ryfsl81
HY1eKY5/rQSV2MjDQySYa4wbhWFPubjOtkfhV3kr8NoQ3o7N3HLk+xqgXkVzWSFd3SChqah25rJ7
T3d9P6ctHgByizlOUNbZJ/jpg/LM+dFDjf3DjtgB7xeoOONzSGEfb/gJxYJjwDfQxv2DkzmHw8AZ
BkkzRXpCG+4+6O0aJAN7fiBC3mYTPOxRfPspmx7a8Oy5WyggStQh0HQAbFLfdjTxDhxB6WRm9JPN
cZCiiCYl5XIUqagL3Ezyk2GDWsY3Gl8jLHABG8qbzudvXI5oH8tMwvsHX0iOpshynwaIjnwv1/zo
M1B/e0OGEM36eXyE2/GjlKjm0qo2HATclynM5/kqBxw602NbOyklWq+6H8se4AWLGHmkBB9KPqwG
JheXuuHNnUEv52W0iitT3oZIWh+HVdHNk8u4LCV3H9uvwOKHfdJI0ys//q4mp5LlQmb3Uu+d7+bT
kWyo/gsVOWrllejb0VbhRtO/aHDnzzo5ZxiDPJDpdhD1JZ6hEnRMINZ4aps592GaBLRGthJod9V1
YIi1gHA905lQOZI7Gkrcix8YrM7gfm9M5dsPQdEJFvL/FDZrOxlCWzpaPMGgwy78qSJyuIaJSa+w
KOByDdYw/zkaugOudKbmBBzblVTrLIS3m4Mevvbkxo0+tj9azM/xXdI6cx3Ob6PiMM5coduVQW5K
1d3SDJe+aLtjB18s0tRZOg2DPyCxuUOluymWxbGTAfoq3M5Q7EBbAslrx+fsPdJlFvntHLihqKck
eqPmlsMBMrRQusTrmHMBWxdYDDETLCXzFwp/iWn/ljXJIAY4vLEmyz+pZA1SzuEleaqT18AkyJzX
njflymyNhDNWiKWy8Sc2D2JhO7KacgvufZu9e0COaMTD2Xpb8uau3Nl90Z4MuoTT5bwHNQCT6syF
Il1P2PzxWoZwRmRkXBaBdEpekqafYVzVHR4ENY3pTP0jBwVshA8n90gpR7IQ0+5s9GEjqmBCTlAF
EPv5eeXVYrYpU5iUAe0qTLQxgqpfmjV4o7erq2sKaCjbBVxmyGdn8DQpe3UPzPlf7I7IKWejq5BQ
g/SSvXULRjqfbNRDCpvVYo6sZLQzKF3pqQJjQF727yKRjOizkgPkINOD4zUIwI+fgVjgFTyLiYSX
YcO1QImkyepZ6WeoZeHq2KHbUJ6aynzxLH9yljkuWh6taJ+s+00ONaZ1Ho2m9g1c79cluu3v7bCW
d70+ItdOI528HhpqUYm5KDXD7caZ/xDn+Nc5j7PwcpQjNUjsQb+42S2Qi/b/z9kN1OfmfLw9qMXy
LIqweswFOk9z0OArRknA7AoBXxiEjKPraISARuDjH1AhWoIb5EFGqEGBBATCsUvpmrm9XnArb/2E
6gAu89oYq7AndG7sgj3eDw4PqS3dESWd/n3MemXxFZPo274khZ5gamWYj4PvgVLSbOsILnALxSWA
mRWghEF9kSe8rYPHnnR7f+9Ul2y4pWaz9TbWg91RJy8LEQNaaXpiX+tD5B4XtGcJIGh8IDurVA6t
0BAZWKbLJpv7jd/dU/OFBbW0tj6kJIX4+JsjjoLE+gD6xIsvgMM7Rzvy/AkCCeI7dgCG1anhVFA7
azbtPOwz4EYnCC0LVJ3Us1TrqFLT22QBfbVr9lcJnbtWcYyUwPl37CekYIftV7aMFk4ZQkLoyAG3
9ANn94nKadyy/3LaqWIq2+qx11uH2P45dhtE1LlcxXeGxi+ys7tW0cf1OUZRnXJGOxnZje4Th0JE
WFoBoC9zmMerVqhy4iTRf2fNqIbBXCsAPZZeFLLASUC1JAgikgC2WowRQCpdWzC8Z6fJBRko/7eo
vi7Pu2U7MMXohphwumf0SP4Vt7B+dKhTzbqyUKHC0O48RL3W/Mms4lc4CI46erCGfXQE22jeNoes
0b51PdUUc3zYWubPtfcC2kCjT6cPYvaYqkuUOXhdGaTJo3sJ4JPSrQhzymdNwBraYuDBLEbbUiwf
HV4C3gMFT34lQj1Eu15uGZV0ZGYy/X5VEJVT2L32AZqtX1nSjtU9FGgFm4kKmD9A5RNEyunJkeDb
nxkzKSh2VMDotWS+R35uY7cHBOoIZZYmWDgNMnOZCJWpH/wllW2HgeUVutwKYSlCi5KWJhXoS+tb
aI8s3i4ASCjsf9r0QyJoE6DQVQ09RN+G8z9YS/njsL/512JgAp1IDFnp8ifLRCTWs5mwg6GPABJ+
dRx3o/xeo7tO4sK8t/IEnrCipy8TV6iustyr7P0w5JvsjMGJApxIaz3PpYHlKdHDntE87O/wPxzH
Im6SR7P4Fe+eeIVAf6S/xyPCgE7OFfBdCC3YllqmmkHHXvmMWAmskFER6QPBPoDnHSFaz0B9VwRu
ViLFMBtR+KiYeaLH7k5RPrvBG5ZoPpLpH2GaZk37rkiaEOXK4KUbLvUQhWPzpyTr1YSbsF+YpcfO
WuuEaoLULEeWsx6w5EgOFSeD2/aE5lvANVwjs23YORHEgDrtfNtPWmCYkqUeKXtfQYY/J//fz61u
ld9SsTrO3p7eREMmUhx+wSHgooFSDe1CrHkhRtijojmBhfmPIvpTC+PlxViu+ni8zkkeJiEMcWLk
/hpeAFu0jtB7OxWt2VL1s9vfikV/DVHv8fT9y4HV4sYHZBMvRCp5Rd99Bi0KjxpjK3sztewotk//
P6eCGTOt3iChrBGhh7CiHdewAm3p70sSt4x76EKBVpNmIoyzdGZFsz+aGC64ougi8mkduCfRwS3U
WRnuxTZdIcW0keHnKcZmk0BjaA/rrBJynhsFbc4g5CvgwPVGsqzUhww5dA/g/KnBN3aYr1znssRd
X5feY6bLs6CfUQGm7gkR+jNEQIJa670U9+0J4zaTpaLK+K0SonHlMZS7nCDlDMUo52sQOtLBzncN
GHD65UYnPEo4qOlGQPA6601TcfWfXa97zJIAiC/k3uZkLWtEtVOf8nIYBpkAzWEggFI0X87j+Q+2
/CX3lpSPGAvJoK68ZjEUnQbH8sI54OI985bRd+7VipfG2ZxIdnHb4Unq/wR+qsQuxUg0Ly//SnEV
2HluIlXJCfLBI4mky9pW9APYv8vhyLu6G+lMt1klIcpg0pspva1xgqKfiVH4fyno+YKs5HkuAJzB
pKWtnFLLg3Vfv5QJF8RaTeEjre4UG1/oW01xYjpsS2CFb6KekP7oSz/rLCYy+2qjBn686i33MzOa
6KjkKV2j1Qi181C7OOSVpsLxNLndzbTxB3k4g0DzTaEeL6Lwt+b0NxTR3J6Fnm6/rJ1q7MOlQGyn
4PNVY+tWbyX6ZuPJa7/14znuAtoE5VJHX7Axqs/jWihMFvKCBaIwxSLbJS7nYuCPz/pBrzClZlmC
vJRDSjewrgVQVXhmacWNBoK5ImG6+3zHZJlZ9sTZRYhOKOxdWGmu5xF0Vby3kT6ateQqI/013yGc
9jXW7IqSDLyVBIIdNoeVLvt/zH/sVbAgSo6W2A5U4zLLbrj3J49pEg/HQkfcKfJAWIISSl1OCZs1
fTZRlLW3x8MD8d3QPxsYBl0kGlfpne3qVFeMVKwP6d9X3jXu4O+51HPXOhFKEUd/Sb7td9+rubmh
4M9wwUN4XYCUCmpPsBSP/RFsK7WdV64SkRH1DNDBW1rtoouXF2srKdjngArMtHyqcQ3v7U7KqRA/
p9z+/MxWDo+u4CKbvMQzjIvKeZztM1OJw5938Qx9us+8iQk3AsN4vk3/fgzGBgCsg5ePP4b0y4LJ
ir3AQ0SH77TXLPknploq5fCc2IlPG2KNL2mq9W+sVMklukME8i7jhVBcJmdQRAi1c6CYznrT21oC
j7Whvop6ufnpxB3Y8PhnNaYmBpfn7dRbXcAg8EwLNpYHQEF9I71kjmo+xdCB6pb0qVLWVdQ+5EIa
3lU+B6AJCQqo3rIy580BNDngyGo4tMZYVYmj1eTvgv7l697bPnN2CbCl2hsvMey2CWxv8Nf14n/r
R4+Rg1oslrVHmw0K1LlpeJ6lkdLEP3hnoxFuFJW4ZAw3iMmwk2dxHcV8TqOuuJbRvzpxFXPSmDZg
eRapiioAnM0Y+7ahUTSj9tl+177XPy/UOPI/SSVeyBiY7WLhaBNwOfj0snOu0Ia4tkMoMItz7lLN
Uus3IfVnwn1qoPVq0ZYxCVUduMXAs3DDZ3ckIWE1UFgP9KNNcO2HeU0DXnonjWYAGe6XNPv3cG4q
BnfresYf9FA/1qDUGlAk4qusQRQ6QEz/3TA6LlxME3/uONY0wInVYNozKgkFUyyoQuBKlvrLWz2u
47STNIkvrpdklt7OlYA6Bd0FZphbyPGQmhhz07fW495jRyVklcrMrO9RmmvMnbP3nJSRBixbWAEb
dIJUGLU6c/WZ/LUA+LXOz8Sypul1UEfVq6ourSp9wLwRr2MJY+NRGL3C/F9JDRqG+NjqHKRbgoBw
EkiMgDw9hk9E6B5ZhqTSYjPCCPxevk3QRbf+Q9xtF07DwY+tPDdtB83yCfmurZzzByd0VRcd3RQX
HNlm+vnEUTP9bGflLgeeaFimE9K0l/zHJh8Y8NomzuD9RriYMbIcAD0FS2Dj2cI5ZR5cTeB3Q7cB
UjwDR7EL88VSWm4cj2IHNxRfSChCDEMIZa+Q5QEIgKc571k8FMBhEH0nE3mMCQTyXNnmIezwTWFl
vrgY0YQI2dQeF2cdyt2cTowMGy43QdQlQCOa6XqPux8IHDSolVtF0mLZTXmYqL2OI3OFkYKgnwu6
XlNv6Z8c0zsDT2flobsBS6RDKeokOHOoIKHWVFB54c3bG46XxAy+NqfWzfVjIsWniGrb57DIcGOo
atc0H/Sj4vgLSmkRoYtsGPdCbib7QaQlfkEuhrGgMxNoZLGaLmJNcGZVs1qJsiFMbLJXgj0+WNwW
OL3mk59Z/XMlo68c+5YLfCSSizXSztxtqk0hLwR2vkptN1cWOLi8cI4UfCn/rqtn0Hc2BtLfTi3t
y7N/V9zC5Hgwbs8j6m2JReZ1HMkrxD4ef1BP17B4RSyC1bk8L5hEsooSC08fd6IHIpQoW2xTe/Rz
vE7IZseV0IW48c5Ns1lAQSkKWC9BDoXEn12qIGU0BXqiwRtITDxFMf9EzNs1f1/TIGz1cw+YmcKW
tWBiUpkrVJIK/Wjjrc2iJHAZXRoMfyGJBnLhAHibHwMJKJtGY0LwUsnB08V/BdscJ0O6LgQM0vST
YwR5PLOtggSgNQ8x+Yqapcl1AI9dcjQwclnodRwPCyqtOYImGCog9Vf9mAq1+WWjxRzjL84qO/Im
GhJD6oxZWEBeCAHflieNQyVUKPExl1wi8u8jSzp4/F7Iv0TJuLEKlp1JwQj8JFqGvGzGwcpo6nop
PrkUhhwtbP5drhigg9ShMBNCEIpPpNj2KDzvBG2aW+6FSEm0icaMVZxacnf+ulYKKLk2PIp3bWJp
icAo2Ri+9Kk/m+BuX+MW7IkjDqdt8s5K3Oy9yD3tlPJlEriY75gGs+639F8PKAz7+5qvKYuEPsMn
pJAzs0SQUxlU4iNWo7djWSLdDtfhYh+tjGMFgndY6hEV/AGLgvoaCF+u5sgr2Ryj2B6D4IfLshch
1Nl3JbBHdTMPp+c7eCDj+0TAq2jcYRdBY1JlX+TOq/Lp+BiDbo6Lco4BS7a+1xw3qkW6lRVfKYAG
VZkkgu2GOx80b+U+ZqJmNomqwCyUdnvvFNppll8np8YkUnM3FlFSTdGc7sk45bKnFVHGx+DDYZHa
eAo5I3S70tPjvr5VGokz7MNg0/P98/6Sl+T8+dHGcoeFXet1Fpxbjnu/0Vx8mwNKR1vZDX3YexS4
DHMpIlU8dtWlqqgpf+hcHQfOikVT7ODfFi32QqGBUrFP4uMLu+1bp/kyji0SvDdrGcwfFwF74aYx
b0WpAp7nkXTRM1kY6+MBtWkI+zdHo5yrx2a1zyj3qxbaeZ1wQFxjQ2WUeGUKfnKdOJvS/xbhVHcO
ys7K5o4P6C5ecTFBfvZUGMYVj02Sk4fn/Tn3xtNadEoZfHWvWl7Dz6EE2ICxKJkexUDNMnXwT1eE
kEf5AVJ7WGhPrSnX0qr5yU+WsgAad0B9nGDVp1zemTgcqopBWkkRFc4bdNUy6Gz1SW4TAc7UGaAD
XO8QRD9qZLH50x7BZ0hYW64GxXYy0PIwTID5k4eTvEyQxI9Sl7VrUfz3DMX1nqJcKHQescrTfdzv
QLxvkS8wdX1ssGTL2JGub29EZ6Jz1TkyJdnR75/V3kWHX02wf2bj142ivsjQ3eMDeaeGFgm28eX2
qg6K5PhhQdB6j91jO+dwU/9CZgpX+8Dt5pbRwQlzQTbBjT/CpcdwcSd11vV6tvCc0j3a3PeNEuK0
87adDhr7Gb1+8roQLJdiqTD5ZdPcFIDDUWXfx430kJ+veoyQRIS1lKeE/XXJ80yINGUqxhmcj2jl
kF7rcwoO+KRX4RtBejV3RGtbAqixu17FXwb9a9o0RcN3/UYHAbbBBx7kAmnAKoIIyRpHdU8apyuY
yo0+gFsMhV5JSzjrXw8lT/a06H5OzWmK5kzn1gjNeOIM02YgwMN4O8a4AWB/1FNVmn6SW487s2HZ
wtn3bfYAaam1ogaA0tEjCCgwwvgMYyJmSzhOFe16Jx0F3ZrcWgPuUZ0r9QziMyFPpPT/4lEx+mJ9
7weRafR/08Gna639jGeC28wqOWVAyFgRKHYZ97xp0QVI9P3sC5ffnHI3zdCmjcldeQe5lx1jNvFZ
Dc04e3aZz9QhhD3omn1iTgpqWlGBF37B7NtPxvwlUO8ocy785BpbZ0pBLB+03shNYsLc7GEEpVpP
rdkUjyx9agGx5u1nUTnBDDn/wyjHErf/xxOcaN1uE12IHycMb5aNNwXKMSn4P36TOh83nlMNbM+G
PLg2wKcGWRX7iHtDkyHTDu+vmHLH0HIaR1HHxnYjjPJMAObV2mbwp/ewWIBCl5Q+CJ7bpKbPCHQo
+8X2Et6WnSvtOp2kQQEoIoaoUBbKzQKCY1DS7aNU2LY7y8rNMz7I5Oi6D1fytpCrqxRIZKhvCyC4
MBRBc4bfZJv5lE6cfpn2eWmU5LESUDfHGdBUMQ4bKTPzkNO+h716NwP3wGCpWqeeYxayHhtLU3y0
DSBMPvJFz1wkICCvDS3WivJGtUcn8CLIiJD9ZKxGnGDs9jBMtLIh27qZyRscPItME2hS5ZcS/ZRz
0dq1SNGmKkiQ8+DWCdswVbPy1tAygMEaSdJHhnMfrBmkVu8aiKGYCjBkRr9NZgLBHvaHPi2WTiBj
Of9SjIJjpvFdEnuAg0jzRrFyInZLtqSriX3LNSnS/T8L0J2nONDAT1Sm9mtYImHAedwZHyPT+1P6
QJeRnV9rx5QA8gSYHgMuRev5YXPPHE6d/jEbFQUZTUt3RWh/ckDgxQkLRyRBRcHOcIDjfwyya1qV
s5xWjPI+kKq/dznzyk0AMNYIlyO1GzDVi8ptBfPERb+ViC8sLVGbKr/k3hvJd8SlrH2cZeXghacB
SMlVy/exXDFBDgZD99rkTZV0Dm/5VUkEfVzG9f4n/jZoBWSxfAJ7Oda04G4=
`pragma protect end_protected
