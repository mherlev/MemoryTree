// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:47 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
QaDCIw/rFzxTYprj3/dZD6vI8yW2Srm01vNS7tmcAXUbjM2r1CF2k6Uw+AhQhO/e
7VuhtXw4pPnyw7RtQ2kevLDuHK/gFCCN675Ya/VI1fNzwYVSbUU2mzjU+BAFuqVo
zlqulwU4urSlkJ5+xmuShknog91xJyeepfB7OwkyGuk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 38176)
+WQ7YoERiZgrTo8A5TNMESHMGSJwxy4z26pTfJYbXQFeT4cjXHjKTvqzdrx7unip
grDnN9caLeR6ejYBhe5E+ufXnjEg7tYpfPvhsOxBk7SIGrG1jizZgMEXvzT068Mf
KyBbwULt0pw5w6U0QMVLfI401IFGfJPyTZVX0Fodagnh0rQFH5oXXCiNmsAKctSp
Lc30PC5b1685u2G2RSc5+5Lg2Y9EddXzsdIkrPMYAN5Pi2R0uhGbU71+pg33sQn9
lWY+bfRqVMlYJjx+nNGmRMdggN6Nw4dpIBupl+yqjSSksMZ2igXd0fcgsU2Qtpso
dJ1RYNqujUjQL5otE2ljJNb6fa5Zh8xT73+R7FqImXoKstiHfxewG3AmeTt7iO+L
2hv4vgucjZ4u4mUadLCJieELPOObJgqFIdZ3ySgwTYKChMILzHfatMb6hxe+ijaT
hTpNWj5BDRQgsZJfVg/wDdU4nPwUmxP51iyobTMxht7YqWyjjc7BEYpi7JBKZByg
02z0x7bJyFz9ZYPEXogAqRGISUX4vd7ZHRpkTELQlYZCHUXFWipV3eO/p8F4Bz1Q
ICIZZ1fDWcGPZpIQxed86YMUeiW/ebh2699vpqHMO2KgoQUaJx8BuXEm/KSt1PNJ
XIrq1NeyEgmpkwyWQeZBjxvyxGfR2hGlrbmnxvUDP+lx3xSclrLdshiFpiP1U1Pi
Us4qQBT0qZ7FEpQ03p+qoIb8cMm69XoAUfAznyNITiJVdHkyYg11A8UXvPFAQfEu
qdT8H4fkjpzB48dTUMbjGvYLdJFWHrcI55WD969cuo9CcoPMHQe3aKvyp+fXgDDO
xUDpkiBgWGNNciQ1f5I/xIpLsbneje4vuL2JAOT1gClEOF9Sl8N0jNju2Ca5/DUZ
21PUfvxE+EAogneTTcjGlT8Pz+dkqUkbDD8CMaVLB6DWlzD/OAvfYPd2hPLjk3eK
7JX80AUAAdsfac/kzCXCuB4z8fiQhqBiht6uHTNEVfisZmbLuUBDWym1qy8ojeLn
J42C35qtWAwPbLn0+bgBM6vneWhMHcFJZ59AVNuA2Ag3K8mI2B8RbJcCM54Jvee1
Ogk1rSNbPwgii8O1aIZi8DzE3izoTgbF3e1sBdv4nUYBK3YAhX2tgOntjAvz/NHG
ZQgaVayu4cllJ94fNkqYsWaHulZV6Xx2d/C8J6FhR3hasT3oyj1R+SWigB88LZtZ
UmQav+VH4QWQWggyHf4ntMbMZrz/d7miLMUfX+y5NKzAemPzGU8UkJej1P8pmmND
ZKVwZ7DgofOQaO/Z27BPYkHmIJ4Ks2pwQNHD8N3gjRry7hTma43t+J8oyaX9Qlza
fWZsd/q3r5piKhi/2gY/XJV6oC8hxR5B7yFdbLdzc3WmtO4VuUI5WmyhS+nkNS9F
UE8ez9DLiikwfoIvz7Ot02k6rtds1h7wgHtZpANbNaU+uhc5MscIPmfdkw4gy2Xm
90B9LIPq2BglGKPk43RGCpDmFiulnzVnDBB5i7419V34HDtDGkg84MHcUrQ6Fv33
FtJEDHxDz4BiO/dMGxlflrz8Q8s1c/Z4coPqZ/naYB8sMOBIWr+09tyPKoyXSddP
5H+wkrpIS0VbS07egdpzu/ps89RDqTyXvyHUbyg1gA2LRunNA/EGm/y4HVOx14oH
50kszckJ3bwtXMH/2pH+BGoZCyGtVRmbK0VZPcVafDaelrmSt3YBmis/GlU1QTSO
3mAseu3rftbKDCXzJTaPNj5vcoVqClsk4ZnPUDkdV9wd2+YyecVpQrhhbtB8MD8i
GHYYHVH4L+S/PR4654+MffBAd/+6MlsccgoDVTS+IzCuxzcD3wUbVzjeXhXyovT7
BpfqK3FxFDtnEYWXbuEI3OviOSqWG21V61CXLBPsUIsw39vFHODEAGpOygb9YwL+
LeAB9zAgoW9TZ0ZXDwJSn4RqChN8b9PtsTd3lRMufymDRqYOOGQzzLgC2qrnfBE5
jfZHN7i6oub3edvxDulI9rAswnnKlhA9EeGjANY9GxhQR01/yWOSW8ZCwjBWBdfx
hJQ0SDahtoI6LjpSp5dQbnu8wD4SXXfq+5AunKxHOXFlj7PVgtZxYPZuOMSITjBu
XsjYmnIvDcJVhsFhzMGXXBLc9K8Zt6uKA7n6qzvXRSCNnISnuhKtFhwPeAxA3Y46
Yn7qKAMl0T6dLVsojYcwm9rpX3Ze9BbQF00AasRRmYG+e6PBotCRijLcv+sJEfwj
AoeJjWUK2AFYE/uCpUPKpew8qHEI0l92kq72a8dA1hqoWEfHFlItrHHnBnZW7Sk5
570ieVL9n678S6nq2RACrD4vUk3CS5yPAkVX685IFyJhmawoJTLwo71hTFAan/5p
9l+94XNdb1L/xjL7ZgM37Wl2hden1ltbMkSpsYv/OgZGxg5I91CE/QeZH1x4pfYZ
dSseFEq1L/FzRiRXpK3xW4/tzDAghhxIoF2ZecgCBzJI4e5TTF0UHuiZxSArdV5B
7DkSJM+/lY+Ya1tdoZamLT/D8v1D9MNnuzgEqYFUYy/meI3txXVTNWDNEZA6yu+R
/nROdZsLywMAzRRU4TW+7Yd6sAS1fKzZmgWH2JI+quYu/3DV+5o9YSZDjWUmtYdE
cwXMEMkY23qFoYs+Rm6mAyPjnQx6hZP5ne7a8yMYx3ocETU7P3VbXPaEVG3tSqQ/
zMX9XcM9/mDSxo0NLXfEAqTDDTTOpvzgtXUAZMAfvRKE2KsWSUhKEjSHhksD6qE0
YJCNysqtenllyMixofJeVKLudiVGkYwXTZCg1u6odtIEPkouRI7S5wOqBMTxaxW7
p4wgJjsk/Gg4HWvVZNqOiB7EFKuHZVHOC4pGnyZjrN2hIPPhA3SzSX53vhLiTpsP
SDKiaOfnLTpu6waGOTWd2OPt4kmxm0gaCY6o47FuMDlMh+OoQh8n9WdiIGHW07bZ
whiPpMgItGuSyHzxIrfb7/8rCd23xaT9g66/kNOQne86NI0xIlhT/mLbzwsA/xk8
CEb+hijNZVvwcHS5vXofg6BLEkLlp/BjDU1VPejMpTMlDMx/VuWmTlLnh05v5t/M
LQ4m9LuyFVCbrAsftlkMzNVzhNLVW/D64/53U5HV45uDsmI20a2gYNZ6LkBVaTDs
i9W9Pyl+T+KqzyA2g2WhBegMSVsST4dp6PMh0u3s2CMWOZ7nwWXjM062fjJmGepo
X5kuO9YsaKbgRZLovT7xYmlIqSiyh/5OnKnKNffxnwH3f2VpMnCPI/71BeCtCqKd
L5LIX0BcDvSgkdMVjm0MWgmkfTH66x9jJGAuyHSjKeYWXlTfLWM0yxWMgjQWMNfd
33eFnV+54WJevOPuUZ9YFPX4SeUfwP2dX8bhP8K++S6+thnf1L0G+qQdA5B43nTZ
c2nXd8oedc0xE35FLsnLOZRqgzHi5aoswf/rR5jQF8W3s3X1tlYDunzey7cy40a4
znQFNv1WmNpiTfWMQ50ep6ixzAwtgkiKiE3IpnrmHBKJBlC1RrZ50lxTw5D217Q9
Kvw+dywLt3y2IG8iE9dtURqdbfdJPViQNU1L9Zoadg+8wgRyKfBTCqWuSiCmMCvs
bdUfDCPye4rQ6L6UJhv/N/4JnBOqbpFw8VFQDjgkoEg91ERh4E3Bkch4e7OgxVCh
BfmUVMBxjcAZZTlfH2CQZzAjaaL2lg+oTLsTk0xBsLwlZaiJU+KIcyCAXwhJVREk
1HoWEZHxgL56ycSK+KahFAJoyKXI4uEe/9jflpOBFPQpaasYVnlSEkP7/Ra4xJXl
t+HwqC925mbQVxidyc5DEKFllxKe1mMxx0pbKuAuPKZSlYg4AKdDc6UCWn79mG7f
tUMkrgi3nIXybcIAZ3JYWhCxw1MNwxg6bk0PwweHgyZgaeNuYlJ0tH4VWbAa3Hv2
Kkk0yh9ldNB/DyEC+Nsl6P5ablXdaN9OWE3LAnSToPdhfo0p9wU60LPJ5qE1mOma
q7aihpyJQXnZSIourmud8uXiosco3uIMX8EN96tpHFpW8ZyUtGemrjgZgCJBy917
UahfUu4ga1v3Biukc0kiyTwj9xHHGQ6CqwrOGrjz5/2TVysoOAXKZ6WoLnF+r37B
07T1mv9kfY2inKpHMePVKSRBl2d8yCwtGWii0LVMKkOLrJQVVEqGYVlT+1pxfAmP
NvS2KfKZFod0GHYYSt1XM1s6/p7vIBUxUAIRj+2eu0yPPNwPC314mAO5VfvSKvnp
9tcafK4WvJcXjMOj/WCBarrOMPbfRLZ/GkBI/rL5t+fdTugbJq5sZ2gb3qYD9/hj
xzR5y/UJhs6306jj8Rw8oexmr6xJGAz91wS7bjECoCb9fEf9XTzYbIGtI9SttksA
Y6r5/sT+Sw2szuc7Ffhwf4b7SavJw3c0S1Pm+D1idJz1QIwByG7h2a0ROV4UR1a6
8Ak8mrMsvBuDbrYXO7xQ1WNFokmHLI15ahDKhXHcNTIaZEe7eAg7+ekBWJjUxJKG
RonHxcxlyDBodtJbUUCOqLSMaqUXsZmmDtzSi2O1NQrKIqKTTTLJFstcFFmbySDY
h9PxQqUAnWo9LXzPUoENuqjJuwxY1f4U36+5LkEieBUGvbZuFJFSCc/VSLYh1/oQ
QNcHfaFv3d0lzb7O7t5xNdk9lZoOU/5yicz4KhRI9CHZPYSm6ySz9DYBgnTr0QSB
anvoWIg0KuX/XdWRpdLv8tI9zi3qgGut6HIiAojxLU4IJ+mZ1zSOYTMdBtjXsaVj
YJxy9flMh1xwHuj4rjgzvoZZlW4U8IRPLhxUhnNJU9+KAjdvWzUMFFequ5WGzyBG
HM/kxKmp8yZut36Flpru3ebdpNWu+1SNAROEb4A/kjzBXIRDIWzXmVk8i8PQwQOg
DhqaPmLp2NSCwgfInppz27+uxObQLF0JNS9j1HPHytd9iC9nrCSToyHOfakkkEzn
Qon5HJ1MGsLwmFu3wlLyM/HuuCBYBmU0LYkWMFlkdLUnSt4IT7N6XAnjdGqdf9Rk
8QZgbhnkhMlnlC+Pu+saeHV6hA9Qs4nUnFRtaubdIuWy5WTnjCmYYUBhHm+B33YJ
CLT+7M7Sq0JTgJwLByQ2g/pXjkVDETx9Q2tYdWny3wMLc7w21UsntQHpD8JoaL+h
WG7QUz/mYHMj9QyfQf34xnJ3YRXT09H5s81dXyECifUJvOjVCVb2hT6K1rMjXLkL
4WRZyRHUvP9MzLG+6nYjapy7P18PCcFgZL3lIheGO2+vA1JMnwH/y1o+tUDcTpZy
rk8yWTdZPzWVVjAFmQ02jHVHBH4JhhejiPyRDiN9b4BAMGuyMw0vpPUk+w6qNfuo
2RFSTCHKF4F03WnjDyH68/kgvxNgMSMggJ9OTAGNtQ/vqaVWANDWACEi3bn6ulyK
599AkJpwOjAX4Wn+9wUuZ6Q4eeNOtjAofK6E+RzXZqH5uvwpnSHgfQqBzIANRJBz
bf8iP9Tsy8hAYbPYTMdWCthq6SzSg+l+OilANJTlj6sdf2+lp4KVw3LQVFRnP9q2
wxiYLicTUKth5HDu3EvpZ7tnPvSIQa1k2ha5nxA1fGRBamSXl4C65Cfc4oZGJ5Rb
EYkjlR1ZaVjPjJlfxL0jVjM0f0EnDCu1is/No4mBhvmRzn54FzemquwgqGiLfWPp
9daYRF2TfKgE2KjfwxiQ0tTMGHKzeuc8dvfQHV17CZw/8nBa/Bqv2PLliWhnxFoI
+uLWngcP6/g8peajN/2JhniwdseK3bX7iqIBBXS3yzY++ucBhQCif5PBQ+fh31QA
J3JlXOoKPvt31f33hAioZfmFVZIshDXVDTz4BPChfzp1QVUck+jlv+ARp/mM8SfT
XmprgEOZc4dMWLp67y74fuHNDKz4VqyjukIVw2QEFZe20FU02YSUHIs6yayrELNk
7SO19A61UC/2EVtaB7NI6bHBFeQjUI/Y+KCuwp2D7nUKOltx7C4znIjj/waPQmwd
+e57wZrsli2dN802elLpIrM1QsImdiawa7Ng1bXO9ybG/sD5mahbt8wQ23M3YfKi
kDrkTl/rJh+OSqLNWoLv3qhc9H8KYj/9jbvXdTlXW/blmc7PHT/MEO5448AwiQwh
fs13yZT730DPU6dM1E32AFfTPiY7xoSCO9Fm6thw41U/MVtWzjpuTivzYHZQiVsU
6uHD/DdD8W2+lSi2Pd9obuK8SItzQbb1btl7qz0fbhGW8Y9rJur32Pxh8QQQEXno
pfbX6F3XbFiCq5ZuZGDD5AZIx/9OIpNPMA7fHv8BP62XZGXF4yoGQPh1nZ64e2E/
XwtND/AQHui1UVDWhnaUNFEPSVIYEtZsFq1QESmpQrj/OnBcWWzJGWoxbhpE4PTJ
RE/m4m+GNtjtlxwNHhmZnOd+NzBb2CZ6PzKMZcHJbr3gs0DgoXJIu0RwLBha6dpt
TTEeRLocIoEXkkQHUqSqinCB0OTro5NXAPXJOahY9R4z0VvgZT92/2MjZMWj2pmv
ovVAIYBcSpZfoCPDhjEoGVubmV4bgQuCvLyBMS6zSLevLhVlUzenPOfEBVQU0Z4v
k67pwTQg7F9zZv3wYwIdzlJ8uCbdeLHephzvoo2jUsiE+Z2u4wz/vQ4w9iepJlwk
ypj7zxW1apmebW1ShamRKEq1T2YKyHwpIYzMPDpkVJyQ5SN/K72boGInLYFARwUi
qn2mcVFEbNczxNvxpNig/xnO9IaUg3GVJPrX6hxNrUMTMv9jhhEr89ZlSftdiMbI
JMQ2nXh45xBQIyx9JCHLuURnI7n8Jh80D5kqAnAxhQUPmvnet0K1eFd3A8qo8Pdd
H+l74fGJ5x6GsJW6S7E0d22DjxircorFzXCGaiWwe/l++pet/F4hNV6sNxLjE9ja
sTHkJpJo13EA2bLza7ZWGt7EjClWd38h08PuCz9lUpqNh2MFxfaW4MirFwUBk3ib
64eHar9R5a7eQBmWdNqrAjlQNvhWvemgehOIbI5evpEnVZLVI/qBVT4/J4tNvG39
EUWaMb2LiyCkCn36fwPJ6Gs21+TPt78l9URh/zwpFSjJenoN9QPFLjWKCV4azxFg
Ca4ZFHqCrvJd1zJblbxQMx78OqRRsJ7nolTLE0+n1HLlN48DxGmeo8uCf3Z9AuOb
Zh5f3Qb5rIGAFxsFJ6ba6nXNmcwC0L4T/koSD5xEy4hSqTeMHPUWxsjuxCpdlDnC
Csnpq4YPwGEG7pEEumnPs69nf0uZCSQydmc9AYaiDR9ueTK1nJ4PHuTYxRQgFpnA
raamddxOU4N1SffSu3t+t30PiOuOaIH8z/tt//7woJyyXdRjmKF2+bcgCe2wYUFr
is7g1DQnfdtNeHbbLwBw1meJoQUxRRnt1rTOCKAhbxunI3P/oE4ujYIFBYuoW2xb
dhU07WTNrzCN72P2IEqMVL50Cu9Sr81Lcf70gsHHqYcHihyO/xlN1dPH7yvvWtD1
6Wiptlb0xTnmZgGCzRAwE/oc3BV4PP46RMo6BAleTIV+xJnb9i/RTUXr19f04uEt
v0+86Ba5THD+OSb3b+bNNmqRbCPN++O3K2SMp47rWRFPSFrGOAn2NP8qE+Yj4nKF
R5x7Xw2/pMnPyvMz2cDyxSOUqLqwdwK0a4J0vYVdUELQNX8wPCniGz+qIby1xi69
T6zRrAKI4KHeYrTiTyeuV8+TBfxDJIZBKIoU0a3Ui1psQE0MDA8f9CfC0rySFa6o
5z4glNu7GGFjchGSqf3jPZBpib+V/pb9hh7Tzn/1oWJRiRcd6KZr7UwjRishSRFU
I6nJ1ngxAbStBMnqXFYia5lil5B7lCwkoWzMTBdEqs2A80sODkGQOfkddB1lOni+
e+VEt16Bx+bW9ubgQckqD4aEMa0c3fIS60WIbRmYb5UYjFNAaGYzB9swMjsa0AS1
zi4pqrQI17ltNMlmFBsdbx8wgiXqIgyooemDbAucRnCJrJPtQju6aQRulC2oVUXE
fU46F3lPCGHuUJkHaF3Rm5Nr2hmSqG668/2JLV3K/1CneA2aEujrg73WTBkRiPJx
8RvsU9omE7ZfPqKSwwhw1pMDGqsnXQsqVhNEyyARaa2BDPXn5s4061qGuWITHIur
Sb8WhREbnoUYDwX69ah/g1gTsxK8tAT67kyF11cdlcv0aAm3Ab9yKz0Inf4Ud+HH
ofNl/hFfpjbKa63+ks3F/4IGMoPugSlKVPWZnWQXW04qg8J0PZQtNj25Xn8IGEKi
yWqDaLaqeMDZoEi3x6sQdTvWeom6mK0NrVdVWAUXElyL3QA0CCsN9ijetBBMTa20
BFNXQPTXT/QPaGMHlqVH4kQfNl+Pj3/q6O9PN1127RWKlPTT7T/XTafFDpHXH/mo
qyxZtvGNjYrC18NBVd7CzT1SRNKI/3DdRig8+EzRN1Jv0mPFzR1reKSRx8Y0PrW+
JcFXbmUghjadT4M+WhHocGxO/I0lZhLSQBcxDryIV6+F34MkZpEWEa+pdi8Bd0pM
9ba/RuVKW05OR20ClZJHgbAUgvXgJLqh4yfK5bAH38efXNFaXl0lbNgRPBDR5JpI
4YIHof/FLRP8nN6ie2P45nx1XVarQDbneG5sGr/MMxJ1uG2dwf8gOWdYrtveahtC
mwsaQwGF3panwX3JJAfI/LApk5jxpboeJ58QRD+n/o0JyTSsYvgAY9/xX5rS7VDy
Yj3XmvvTYpk/3n5MaH3Eta0YbN+115tEZEvUnyl4zAFbsA8a+/1Sm9yH45SFqRtA
iPTcDnM0/cuyCMLJjSwI2VmcAwAdB7pMuP+TSh7bS8nr5VwbWmDQyqRt32nHaPAR
MJUXVKj3dAEdN7fWoSNH9gJYWqMHWO6atWFbujU5pFDk5OylhHi2wsCh9ErHcVv7
YhbbUnERynIbnBI4IoI42QP7lJ7PUTSB0U1WRKL6HKxeD818M7VaxMmNtE+9xGdq
OXnw4E8uaP81sKW6xKDJ37eGm2W7WiDzC6B58ddOQ9i9OQCYwvNR0O423cDi34f9
HNvGprB+tK8MrNt9ImCV0v1V3kIFor7BLORswTX1MjYvZqvr9CnSiqrvZ+5dd2wu
HoFdN3l5YG2IENLFoZfzR6Aih81hD4417xyvK+xffvU5c599ugDO1ffG3Afkq3o3
r01bs+uqPCuuUkUbzz02nzpulcCBIq8B+giCu/l3E8DInaFlD7WKe447ZaOY54tG
8rUz99zYVj5A3vxrzQTAfmMbloM3AGfYXGSNRzD9anwBJMX+qndFRkj6mkJxkxAg
AOeXQ+tG2EU+pdj+LhDRsa8xEQw6RmN86Ee2e2uGgTTMj3q9AH/OxCmEUSfcOlla
EvL5BYGggdnh09qNzf0IZzLhhvnKbyHQSlurYnbm66rlg+4kxB6PkclxcdlVBlcE
0BWtuPWpiYtnXG4xKIo0KSMl5RqIKXecU/jrskJ3CuAaOjWxEHNeWTfGZ3WFdgxk
JaD5Yr7mcfNguDg6ebds9T9j+ZdmzMD/lKD4tWtrJBOKIev7pR7GVW4xneD0935O
lUYLlYEfP97dGy1oZjqTwsDI/9tP5x8qcvFGW86ckeR/WuLPGZhIuqu9t2g9rfUH
OurRfTGW9Tay66lBnirMaNKwVjO1jgLFk3yICBhjdYyApfp9MWNLnmIkdVt/zee/
hu9LDGe3F3GUm2963txKFSwGcazJY6be0m7cpkDLKshP/VM0e2ef+wbU7vMVPrIL
zrVTOr7XLii9mOlpjNNr95ifm+3fppdSjWuXTL81bEP335P2T8WH6VReu2ThZezw
kZB06S3I7ox0/3kPYEKJ21/XiqeMBgCwKtAEXwsdGRWsqyY0TacT8tiYXyORtoRd
3M3FyD4Y3FimfzN3/Ye+vAmMGVfSiPdpFM1ZT8VrVjpzXOyFSx/menGmSVVuzQMA
5WildKS7M7Fl+uYS+VnRjPFt6AWxi/xPCJggj4cACCAGfMsBCqYxtONSH7ybhVtV
dJ+7x+9PPB4aaFaHwUTRjl+iEuPSn1FADNlq/wbnYa36CW0aWNDw3qie1SpnqsIy
Pt0h40em6gbtZZVtVnfRotDSTdoiiFwJj5cCWxE1vYh0QovZEdsia4W6mzSldcpS
4UzjVX6ACQvcEVQCqm//A2rl1vER6Gn6HtJJQQb3trQeBnjRuNVGs3o207dVYnEQ
PQHJ+Q4Ckyk3xObf6Kn9J7OO7HJU3SfU6zuRBVFdPHjm9qcotCnW0e++w7916BpP
/k6L6CLVoPRz2lzZNGgo1RuEi7Qg4Ohq6ptaplPYGChFDitRuy9bmy4ciVnSn4YZ
XhFZLHBqzBSn5E8zHiR1fZRBqUs29VuFWA4ZpHmuOqFzFQ0KN8Fu3SBIfNsa9f8C
AERQmwk5oUz41HRJVdtehlpQrNrQ91mNHpEWQP+bQFrVr63GxqKAvzLDhI4bDW21
32o+SaLBGutEX2BB3Z3kjN725As7CVmC48ux5Q1ejvxGUyOYWVm4AwrtPfeg1xYD
3V1PtbhlU9/oRivSF7GxEry2jd45DW3+4mi7hanvLWGKW3OUO9ggWilHqMbjLC4U
QCka9k5/z33KpVdGtoBRvySbPlbcjcOsjoX+11OifHBRMY6APV3oStFioLjZ46Yy
SKW5gbqMgejxX9JVkm3Jpm0Qs6vASHgrXq5IswEbBJxbMSSQLxL8KP4I6YB6/UMM
lYObDQDYjFUYuhxqCXXnSXjyR85XxOSSHvTT0tfSYFlMMcW/d6sqRX1FUxalXRdx
Q672ktPW724pZGZPtZx0q4h1tb6v44yoiZ+IS12nzBVawxv8yFtrGhIEG7j08ECl
jVVwAyvNmx9ui0TX8AxMQy4iG3RjYc96HUG8GgDH88hUmjnhRePXTkekTGdBizAG
aog0Npw4o1h/4ph68ZnYjiAV3qc8ZoMELncP2ZMcyenNwceAqqTDyqzHegaEjx64
HSg55IDgd9lThqxeuyZvAeNlWcXYwy6yZYayuwpD3BmxeuoAMwTDT88oJmH323g4
wVLsSQpp1n6wrdfUT96BBkikL1pmB6Cb+fd68xh9wS8RL6dbreV6ej4aGsaBHZGI
ulhZgrCyMhlW9g4DPl1aB7SwEg6JfUGthNSfA4/5sx+G0kDxbVeYE9WDxSnO/XfK
Bdzp0Sh+BlM2UIixjzamvUySkzVObbx6T/IFPdSEv4eN3Q+wOkz2eEtJGu8aLJp5
eZusu9RMdi8urCzBrXu9/EId2Y0AV/hpF7nrUHphkk1O+vNj6NX4U+uoqjlH3RIS
AIKQisQnkhzrhcQPubBYxw3jfMgN6jtog6JgVt31b3xvZySIkbETvES6dgmsVBYU
SjFPAB8IY51u8HOMnnFOyDDY5faLRGTX5Xkuh5T6tZqkPereJh4NFnoGztKvjSOT
G/NAYFXPldZKCwca0a7QnGGRlYCgvM9liWPyjNVDqbs9eT2m15vO+z+XAdF2XLgl
LwEjElfm7vYtiQSqoLlZg3pvbOA9yWV8zOzo8h1u2hf9blCvJ0N9oorthD9NJHd1
k060RgoG8Hd97KFj3N6evhorsRd+pfM2IXP8280AKg5mFATKco94SpNxvaLTv/K9
vtOdzFB23fOrAeLz2WKx4bYw3GaxOIc+vEAbZE2Xc+nSVg8XrSbSGhaVwgC/im67
pt+YeKDwbe2rnfr880LC/NfL7RCzlpf1koVyEdaCnpr+jai6bzsfqYGJU2ip+OK2
xRYohZ+/FbxIUGjQLi3OIgUsLXFcGsh6nrLG6OBQQ1MQwvZwopZ5DV3X2lcscZBH
TEGT6FmhIm+gL4fCORp4S0onmoHf4R0rJjnU7O3no/Pjzj8Tn4UBVD0UBxTj5iKd
1pGiUxT9+/78IYQu1wj5gWqNouayzeCk6JuSwZgqWib5dr8U7tOs6BnZHOvNw5RE
5o/yA56Okd5V9Tlzn6OY/4FKsIxu8S9n1emYLDWxsoAzsnpTgOiJyNH8UjKRgZyT
8dlZGRvohPqz4gYsuS06XiA05TJpCk4onMtZ3zLa1wReFPDar7jq6rwA9HgTujNy
QSLxdDd2WHFjCNFBEfT6rrgwbsi91mk2qpjQlpjcbIYqzTIbN7R9cEioTnmJHbTn
YCdiZUjdaFrej6N9cKo3j35dimJvecxyS3zTTqT80vEPfhEe49cr22uz9UQ6WHHo
6JLRwm49wrZ0JxPmbruSq5zX4jgIc4eiGzNMieWWIka1jNtB+Y+nXbrUW81bRC4U
LgghrBRF+I0paJV84DsYl+Jkj6fRCPP9Rkbuf7cbXi2JqVnzeAF9yZA+8q2VXTwF
RUd7qECSD/Sq1Gppe0lwXBoSDGqgcWCMIlyfl8j+35fbByx4b+iExcJCBdPjDjXJ
xPImgVRrsH3K2+RktPdv7M+PKRa0ibc0Gtsx6JGuRgtHrNhYvTbityQzHH7DsUis
gL0E4xcAdShGsYD1rskoTxqzMaeLGOCiwwuiEJitYreuyMYf6c5R0YVkTDSipyoz
74f70OgQnfcAhGWZj0MOvtfmZ/5gj3Abpef6kwmNe8uGk60SGikCYl/jb3sG39GE
YzRVKz361ZcFLMtRekR6wdnz1TW6zwE21Rozi3mytL/zRnQKHdV9xUVmv+j3nWaL
nsuvLHJPIs1r1nyTMsk4SOFEW6U3+BIwH0FIIzK+C2gVd1SN3AQ7LnZ/nOmprPP/
2fJEQk/zvw+EbEO7xC8+y6QiISq1koWa5ptEb7tgcmeLXCq1RVP7+WrAvvMQF4C+
lrn13M45yGBx4dQRjHYo/E16dDviMkDfsXXmyeEaacSYgcvh+EKTmlaMFiw4Y2sb
0rsNcw1vsji9I3C/6fCMTpa7GgJGTWMr9BUEcPgHY0Eqoni+Vi3AlOin2DuWsjvn
xvTVqNpp28b1Lq8SbYozpyjqLfJ00T+dR0nArLiOmu5D4gQEF9ME1QcCeLgwgQ78
w5bwOGXvOQFGS53yqmXjq10J2/x5Err+rhKFXHn4SM2uWGInuDqOSZGF9VTP2L1w
AREqPC5wk4lQoyGfcntaPge9gUWObqmCu5pjkf+5y+cdUQOf4qiFRSFjXdW9Wt4K
fb6JElp1Av6rXr9Z9bvqp79yRlcFWqSga46m9DAwX1DUBbGcpvZ+BlGxuVcyDIdG
l1i1C4VjSlSBXvNFflTnOlSU+xS3S+eO6KdMZYTG8L9BALRZVALfOy/zoi57UQf4
zbE/lbdnFT318aSFxgqzSjTdBp0yS/PLz/Tb9ptHhUHlz0Kj4qYn6Bt6gYR9r5VL
j1o5imqS1792H6kfrrHKbvFKwpzoEljLwyaFbmCWtqWUOnMmmf6ykC9U8+OGKEXt
Zo62fyk05OaO0z33L3Y4gp2Am4dTf/OeJwGGKyaNbn0AzbMz26wgkq0JDKOizJL/
XMDHws36pkBVCQ+DJMRQ8mviXezP2kyepwp7u5z7+uJYjYdG9VzeyJEaFkRfjRVm
qcrMWpYZCB5ZiYE2gHlrN3HKflggvtdwZGGu/oRbjcXXilWWbJDD29vM/axxPrIF
QcYirhbOmq6AubMmH/2RVU+h6W7ZkO1/etXrMegRkK1IxhCVrp6DdonZkT8qTJDq
fq9uiVpIW8pLgpR12DAQ4LBMAKA4GYHXIQlo5K19sAsCcEIqm7o+McAq8AZtLv/M
hF0snk/RMdwmZOaWFvV9yzPbe8/e0IBBjJ3EKWO94V06Fl6S0BAwKSDZwseB3Ijz
Bh6BZUwTPAcEUc+jT84SYqiQXl70vl46BnE4zVZcnxNp9Ka6gCVZ2bAq0NwA1plz
7mvKiiN98JR/0MLxRoa8puxZy80BfyGjaJ1eETcmxiKin+w//CkCNLddZXGTE/vi
bjvzZbjV4Js0KDAng8ZrDviv8ZXEIqa5JuILcQ8IFCVgjZt3Vcw9jtLnntyN5A2w
LSB5rz8Mlx4U275RSNSKD8PtYWfchDmWNUWYY2keHDloBZQbqD+75CMvMVGA1qMt
UjUf6+AzVDZU0KA81T8vi2Ja3JB9jGsh6FOJVuYIAJb0AcQpofxoFj+IQ0YoGaiz
gR1VgAHlOMIdByFU9BtupW+C75396JR3ZEFStEs6Th2ZlFZf85YoJ/Od4G2aYCsj
Lsz80Ajl+udPFrPbUVAHxZoTK+YuRu1/yL1JFmpi7E47lt79suySFlv+Fl3pKFSu
pv251zC+Rbce1DPQmcyizIITDDcrkbLObln/ZYRe9WnzyGrNYQVfTQq5weghGU1A
LdnuduD9+tBWz2kz0nrmPVVmoQfJIThfQJIbXC15PFPWlPsU2oOq9WaMvVO8NB/o
MOqxQP4/tKvqb5bvgVJek8Mc6A88vM9mcp7p/h9wynPDX4WTLHTWk3HbzPW6KUG5
02sJjAIcD9luePIrFliwFUPPNZibxvUZ7ktez2bj07nGl1v4Mgw06KhtWcwgziHk
Wc2q/zfuh6i7jVluLQPVelPB7+bBwnid0kuICxjG17QXW5BXfv1fe7y1RGrFwJB5
7cXnCBYm5rd1S0bG9XJJEJMLoEkuPbxFKMH76trTxQHmmJA+UN7I7RoYZEkdK4xY
aIXlDqokXw/NDsRJmKTkPBsbvSdiwHy4nA7D40iUMPIWfwzfaIO6HeborzQvbQnV
RYZ9gFiSJciz0BO8IYxtWDP0BY347K17gURpnX2MkQAx8tJ8HGJt1k8u8eY+EBGg
HxE8leszeywAFL0+zAX2LPxy3vQ5F0kEB9epDBmuY/SUBy+u7NEAd5pUqYEU19t7
qPzYtzo/+GWywUMk4L40lYBikCFhgH8awbdmpiiFI8A7t5h/LYo3HPhyifUkmwMF
arsTK2aqSbyC9p7/dG3MnpoqdjxYxEqpR2M+dJer4HSQHSkr6Cn/xoFs/XFF7FhZ
vEAtg6cg1Jv+vXjCWCCk8zVwOgHbiHy0YliQ9R04VQL+pJO3zpJ/Q9Z9uDVUyxcH
9WsCTANO8ljJ1Hs7OKSSb4U7MKh1l/3OvpdUrA2xTxcaNDr+c8gAD6Ul9MmPU2RU
DJT7bGa48AZeMKN3XghwLL3t0Dbqxfod19seE0ab+u8tHTLtEriBH0B8CmOKI5zH
iMWwaggyKKLZauFpJeixdabBJ9ObGGY/XNstlX0gYjip4QJJCjmzI2yNpMarMNvr
mOYzij6/pj2Htmj9qf+/BxjCI3PlW6on7s59Cq9AbdwY0O+VUHEFLyBs7Ug3UJJ3
TGO/ZnroyayDBk2Jytmma0dHWdVdiCyRBDtu6qaNvtZL0yIl4+QacUEbjSqalo5D
Tu+DGNpUR+pzs37AwUlBCwxU7B79Y8Y5eFtcn02w50FqqmoA7jXZYToNjAYBtSgo
lgP6KNvzUp9wWGL/3c3gjdNVpQXROO3jLPl0AgsLfdYM/wTdKz9LAkDWsR6lIRUY
ZjIwpU7+XAg9PgK//AOjXNE9b+6cpAHsrCLm79y3le/1YEMovRwFNHOfqn9XOkSD
Q/svnqXsTsVDs57MwpVmxERzHsNpERSUCs4Jqlfa2I0fPCv+jRG0SjBU7mlZK7lz
NYWpNpdWAkclDnNCTEuIQOjqcH/foUGlmfMhL0U3ZctVq1ifBLunyF/fr3ebQHYp
uPLIk6FTlyHKfgPIMWf+vcRJYbTFfaXJFrWUkE5PXRciLNtRLuHPMyvJFDuVnnrP
QLPIIq73d7eDalJOVSwtYK6qo8rIXeaG5cv0hqOImOoQ5AFupkrSihSnSSleWROu
s4lPDAEqCgQSdK6H9C/j5nsLslGtxgNJQ1GJCVLjTDmSOGuZfhwgj4D8KaI159ho
qrhiDRVlNIV1KyXuBDSxS6acf1O3CiCYjr4VXe4o8NKg4egRNr+ka2v4CSPfXsIK
P6L5T0NGXrSstQvh7X5y4Xcu3h4MKHwNKUCW7IBWwUEm62/YSU9JFAeSrVQoBkv8
QDwNdScaU4izREqSlNZGE4PUIhsUbojCHmj38nrDChMQksjdZ7ESuBFibMxQKOJe
BYwjyYlchGWjKEvqeub3aJJbhz1Yg8shzgeheYUy9L28NA4yS7un/U/lk9l0UiHr
gctgNFq0HNKP+H5RDKF1KwadJRQbwhHfrJtu0VzLpf92lSnragg/NUJdlkHwv16m
2VpAi8WSdVT5ik4aEbfzG1gH2PypaWDbJbmpNudccq/Ekl1/OLSsTxFyDFs/lF/n
HgRx81gnMfk8VzvfUFWxeHGP2m2tF8bf7w8AakO1tSEPaKRDSf2czGcrE6LZu7PP
/b4zn7ynbO1GjODo3g+dLrWKhIABVVOExpXgrEO4DHJg42L8SDfa2hvbBUADtkEd
SqryJcEGM40tmZen1UHPMMK37o+Y4Itl+PyeRVDvK8+IWoJi09H8lplbe1MDx26Z
hKJo8pK7FSnnA2OeSlwPsfW5Q7aQPiIok8QsHJltLernKPoPPU8vj4qHZ62x5J3X
QCp1Bs4qkGSGLhGTcN1SP3F9BirIeuE+Ic2qTfhSjk6HWn6x+HqbpFY13sXFZ0RV
YQX+xAM7LB2qH+jodD06wC353VQr3tbPBLlW/5Pj5n0gcVEBObJIIyku3osb5Msp
b05jPy6LBBDmgTTG+4lTMJOXsXMJznDjHEDGIZsYWwzMPJDZrHJShzBayUB+bPRQ
KDUnMVtkXY294TNlpnoqTUFntpDvtEIr8ItpdxMAXKFE70qQfbs6mtog0gLudKTP
U+7ERJIa7/shVqDhA/hABpcoJbdqAv8bpT0HO+HEYBmvp9vvN/HWwTMJVtAuDKhx
8AZ8ApC15ozFczBCDJW2QYJPtNrYA/KCTvGxAgwZb/u6LJ2YLly2tnhAfBepPRbs
/O07ukloNGNizmvpga9B8l67I2ekDE8Fl++ZpR4rlqepQUkEslUZTlCHKq8vAzq0
LHUHLnR7MJYEnV6DP4Q3lrTZRt+mR6Ax69k/IqjW0uHb1wdlOPIGEUy8IhAvcLjQ
rtxB3h3dWns7I9fL+2LW7Owfal4X5j5fPgbFMdxeFfzqp2pX5zeXScnr1MwPSULF
UlhklA+fUTy6k99Jq4JSni+MP+/D5/DV7PWV1SpOuKewLWS9l1b1FKAcFUhyxY11
QUe7+Vzxh+x3bmKvvxuABCseMWTHEPEK72ArfEKjrvRgQH6nojd2JsrwJ1Qaek1L
Aaqu2mKu8om4f9CTTSeIs4x8zXTZBAlj9+4N0qxFGVLZ/krqxD1OgkTMkyTljX4R
5GUtOKC+giaSbZEgkvPoU0hPlZEgIKlCUYJ5bEewpTE0UdJbBYKACUGrAad5lczX
iNiIsuf2SLpwaIGrIClkiWJL6opd/mLJjZ8klrLBlDE8c0fb6HRYxSU/rSqDRkT1
1diAMreLUJ59u1iZCs14fxxX44ojcVjWcdtzQ/xxYxfmuZTsoEEQ8Mj2xT+wtYBZ
xNbQhKGoFoePn3saP05mwS7nM3gzb6HhlZ4pRWch5GQcOZEtzcvWlQsJThImONU2
1/HxhvxVmDHvv0c+44ah4Dja7mQqtivvZZ/Q1f+1hRiomJsBblcydMtzInc2cdEf
pINhdZ9DvcSDigminWtL6UVwN9qQ7FJfKi32pG20+22lk+SQK37dCi3RMbX8z9QG
PcsCzfLihnrZrc2ghPbWCNncW/x+MKz7HmPCzapFCgBcXVhMJD8Hmbl6eLbdrjY3
4c5NttKRh+wRfTTYDsDDU2Zfdyx1z0SEaQk4qMpnnJz/giv8vO1G1zTufEQ6zdgJ
7ED8ttIJa1Ft0tBGRgN9lJku26mvW8AkziOT0GsdccgJiTZ0mHNqYrcvRgPfuIZU
ljdrjSB79atk9wMJXxgyczXFV/9kVEXr7kRuU1zZuYTF4MOHo8tZ40pqv/z3yezn
yjODczEQno+ZNgp0ItD6tBRZvxc6kpTEzH12hC30D0CKP2aNPoFToB09S+cxpF4N
gP+gk5cvm19JnsJDiUb3KWBRrUanqmdIDkGEgp+SAujqufPYA60UHUl5VBov61pN
9KSEbe5yVM48FVP611cL1JOTj2dTmYT/PtfqGqm4didfe/CNnv6wOTryjzY8A4Yk
Y+RcWWoRjQmPRwFqBHsBPGuBTL+7ig8x+wV0C03gWJx5J4mbRQXj4ZJMQOW3x2Zp
VIgEHaWRzIZN03/YmEwIDCcsR58V14GW1AIJUunZ2pm0Ciks9cg0U115ZrvntDpQ
P+AmbTg9dQ2tPapf0I7FW9znb7U3QEH+ZBuA1GZH7YaJMCumcdAJWuRc/ibMYjdU
taG/9KW3zrB2j8iXXEUz9DlT98mpM3Wijn8BntzxQRHAOy3MPH9XYhmyG73t91Wc
7L6givBjMRd0OykXYR8V/vUjcAcXalyZXo0xZ/H8yve+YaiLr/NHu9w09QCXw9kG
V22roWHUFkSRDr7NIo4HzPcnyCN66gKb+g3bPJYmfTknzSXgi5opqucn0fNy1ejK
v768PL75QQE6zyUkt92lAb4WSRtJCr1xTOOGmu4i0/LALVZ4h08V3/cND6zEV/x6
y0ykkGTPchoyAIWQ250iNMicEAFiUqCCHFyfcKlCMwg3ofkjNTujmvMO4bxVWcU5
ZcXdTlqWM5RqJTaP7wlTjkYKu7XkVHMzldH2C9BmNfNdhbe+lxkAEJ1X93iUEYq6
bUpKih/rLlzPH4U69L6H8YBwzSUiqsYH6jvsEiCEE8QDFc7cmqFp6N06EWNdLWG/
nxBxmn4WNQFzvUKala+dTCbK8DfhEVgqwjBbVPiA843kBpaJVIKvphg8k5CyVjdi
g5yogZdI0egEfsDKtmbagacLDd1t7xtoiSPyT5/rlcZx49qZdMplsgIjjTd4af9C
vuY+jin7G6cZowhi3/Rn2/maK2oQsUeif+VcG6soWwcnD0L6/OGjbTEdCDKD7YJo
DyILNWiL4H0i5Zsuu1kochdkOglUomdiwC7PU1s8oRPnUIuzRtdTY9excVEqlLjm
Kl5U3btWdPIQ3o8BlK+j4LNI+o9masnghTFOgTD4gEOd7QGg81IYmZMdFTBaMVIT
I/OBhxZF/F1A9zM3yGezrCyOkdiYfr5C88FO05cNkRq3bdOR5PHnNG/S2KS9IpGq
vFYZXCMCJoQp02GBlg5CpfFGfu92D+MjIwcm6UGRXF3gnQESsseQcBKrxgK2kTNF
huv3hAL3LbGLO7qAezadYXVrdBc01T5n00WzblsNKc81IQpEWlQMJyZjPpaoj+gK
WCR338/Vq0Olbujl8w6IigBaeZdKA5fLFQ8hVNpZ0PJqcxOyCrbUdT+9R+QLSkow
bQn5RadUYbVgvS5LZ/Y85g5MronldA8IJFiMicK92XqepPLJh7TbG2x8+D+4SO3q
BIjZSW9iKh4cNrkRYO+2npbrfLUIgL0PmDtisKe0oQe7+uJpMHW1/XuLKXBM1w3B
lwfMVKBTjpjOom+PJ378p431+HhcRTsCLXowUM6ISJ1iLERdTrmLaHabCF0Qi6wr
URxjggWRMKd0LdoKdiOYOKXfL8dLHGm0cPzuUwUTBKQBi5U1g+GhU4X7pU1J7ppn
JRipTni31Uq+SBDnKa3HncNjlCyonqucFTmrajZqP/pQaE+/i/C6Bo+ZBTa0DL6O
qwFPVEmPqgx0+3iTFS8ckJcQTuB9TUKB0uj5FbuIojpJ/pK/hTibyhWYiqLAS78S
kJqYn5cUpM4kVMuI1SVL6VN2r3Gg5x7kQDES5AWJMEZ3FWvZ/aLBNn2eRFoJL1NP
1RzVhRYhK21bGRSA09IkKlawklkBeNlrFz0meMzDGE90UYTArr4OXk2URDrsfjb3
mdFbDN9sy7XjJjgLBHHDMTHD6vlWxkp9MOqnIYFUvwD6J3eFkCwD2rmbmO3vVEhN
LiwMIANoVjynhVhgGC5Hl/+65JMA8o65se7Bfz8JTHJLbYA0BPqTjbctStQdRp9W
zG0xEFpXeUcU5QQQO3R4NcWWH+5Db/OYFHUNsL+H+NUnNmhafXaF6okJCVuaX81l
/5StMxMzewYNSnoY1AjjP6zYGxYx5F0w+n+L3qXgq3j/8ssXi9F6Vi/lO9pk09mv
N/6suKMAaV+vuSupbxHPghmWTiq6Ub/G7v1NGIs4XAxRapZjBMznS8sXGIjA0v8s
gm7Q5bipl8LZN+xU0Z5Nt4Ao8Mq/GhN+dDAWOfd/1pKdUxDrT2PQ2KIjpAnNFeDh
5kxHbiWpIaXdo6dlCifIo3abPG9Mag5I/qe1uNKCpKYucHOiX5QpARQrhF37J4IF
+SVes0NLLFzo3x9+Ybjg1jkDBDiGMpQlrR3Wrd3qxg8/JMpsDeUGZKCawBgoLTai
hAU6+n2X7s5sbgANgV5Q+S4Pik6Mw41UnMFD9L3CDy2JibPk5fwIC51nDE0tpc32
fMhn7qCP8/KL4c+UWkIAZT8O6dEwAITdwBRgYJfqdZR0c1udQftO5JVdT7hL0bpG
0GXz8Ato3Lms3Xoo7ZsUWbskMtBID9cfF9Hr8/tUuFrBmDrAwYMiXGJow9zJv8zh
yJTuzsiq/II+blbh0vUFqJKhMCM6CZEi4DsP8BTdbcN+zlsezj28A31CtgO1GpH+
X3Ye2hUb6lnmuEEKysFmfCyxQfe/GVMy3q+J8vflAvrfp+7mC60liweUdBtyHJQ9
c9Pxqe1YylpLsnhBvxfXhKnOZQzF7UgNoXE0TAIbxwTzAa6pN+PlWs4W/CWj3GOG
5rtCxH7wMtwTpqbKn8OMW3v5U4VUk+bfJsKnEZF5Vnfef+dQsJew43zsJmH+nP48
dYpy2/lTAi5Li0gFI+CdYQnLhHgQmnZymac8xqIwrNZrPCPfRl0SAPb53KPumbvX
TzzfBTnqkxD4Ju+zcepGY1OOMh9PVKcQyfMO0jPKWLGtR3tosP2GW7huBgE13hL/
klKqWep4yJij58ir9xil1G3tEmwv7Rv5mOW5C7j0JIWOiMHZvskZGYQRcrN+cuc4
hu13C0WjRJ1IdIiFhHORlE4Kh97VQQCCjJhBqwOtmP+NtyLqx7Jr4k03U91/RBYj
4bBdDg1hR4xZb1SPIQrNH9ALqQA2KEIeGoC99CGreSsGhGqqBabCLVmWPmh4fog6
3KQ2CQmLR20r0CkFW1LGpPWG06qVsiXdqoqH9a4DU4p/pFgsMsNKgG9vYWMzdQzM
hxrvSuepflmnqgjwg22EawfQMXU8vRmahbgS7xo7VnOeDlszzgrLwBKRaTrVLyD4
HTXiI9rHsUlgiZ8t4zG3qJTOT6bOYHJo/B4mYMM4Y2fANmRXk6t9/NY943aTrFuk
A1ZZeoe9xckB5+vERFp7vaMuAXR9T/LT7mT+n1BEEhSTZnHndrFRvy+1Owru38kB
mYBGfYkHmpzdkoBwS9cTPFwf/CeL1cDhylb9fxpGfoL4gIoOX/zjw+a4BpQBcYRJ
5MZRjMt06DkMnR5K9IgLGRhRnwqNHzdjbjCkSS0iReQMVRMh2YC6zdp+43njD3g1
xQ0w/bPuKObQ49lsaOJ/jj3jiuG5xY/OzmgkBntIS2QTeHO+8/9carMhho0yXeDF
iUuZ1cWzM6GxD7C58UMJ9MD4S6R/gusgl+TdQvZBXxN6Up6HomuS/7sb3vTpoi7U
ESZL+tVjsrY8eM4p9s4Mu7ZTCNa/w9ooCznd0kRNAPkhjbiF2Es24x0kBWxWtm+5
zY3JYHAWMQ8u9fpALRw/6fjB8Vsv62F3FhHJli9Zx1coORkP0ZwN6HI/SfblfJ+Y
kv7T0H9lBMBrAbD5IsPR4x0azvT5rldiEbMlLVbLz8Vzp6XfyM9n4FrHUEaCpB9R
LfA4I5/1ROoanXvUz9zDEv12vJpijRUXLxZ92rLNwfAER7BcDBuapa9IZp+6a+QX
85fvXV676yJv3YVWIkc3CZ+MCcPaZ7hbnGSuNA7+wHuMuyecLsl+PlKDjYUGYW2g
JBtsXkZjBBQtt/K0rQi56TyBqw7g/aRf+xrCCGxjA3dR+CkNMUIJoibJFlASXgBj
3CQtaRpI1Pw6bInUUpl7iT+W/qUoctc0fazv5R0J0jeY9NmUPr8sVOkyKc7UPx66
Z1ehpVqVYXdjVbmLM1+4puQl8cIMlxQDQxm19u2n3ph6XuRHzc03rEloBbZFc4om
g7E7GTWZIiPj8TMc2yIGIrR5HLpzTnznLpxrhE6StSceo00/pxkg4dbJ+0Fe3p1x
7qoplQ54sQbn4YEBNMX/dtXZ2e/yvpOEQaPVmgmBRjIyVhTmhINSD2eU0gay2zj2
5J580+OjwHqSlYt91sk9Cz7tsgwskaQ+0+QzIDoj2mGlJ23uNH4UTCbHRwBlU741
WhvpI/OXKF4wV3z3b0UkjWHq9FHcYw5sKFjWrbsLb3eyPcV0nEZVKwuP2Motu0mG
0MN3LIQphhuGPrRUHcurWl24V6GXY7p+Zfp2PU6cyml9GEcMh9C//H4KkarFLGSz
Nm5kq/BFoo+pDMXP5akz8Azzn4m58l6htJGJz7/1Nd/snkzM/PDzi8pXI5LPLaSK
TN62tiBgyF4n3l3lr2pRq0QXK8cigq2F1U3ixSC7d+C5XP0vbNN2LHO4WyemnZWL
Ma03hcnKPUziCMTv16Zf0nUKFWifzzXkQSVomx6P5+SamWFBnVKEPPmZAY0aPPEc
0fWzvRSVu6qR6xFSqLsvjbcBqNVAcL3j7Sh8sw33aAZhXsEyMZzV6cdfdDhxf4E7
lCGbewHPLvCWG1XtLkJY7EgGgFtdZs/Q/RKdaFwHyquCTI9WM47qpFrW+VXumNbl
HakZSS9bs0pKsBVzplCyHu8PSR8YPfKMUFpGr+EJcVzUs/a26sJ/cRz2PSUBuKjm
dCbDcfr0t6CtbsRwM/ctB79vaU9gQnCX/m5+nozqa9lnPTHPDqUQ6xNtrwRWFIJn
MFqlgHNzYuSpOd+94Weyjm7MbDzhd+Fs5jnCqGiPKIHfoE5vYwuXBw9hF+U5cVfq
Ohlc50fZYldBUmdiZS0Gbq0DYPOT5EGy2OnK/Jzt+eV7uZ3SFxc1tLXYnraoSM1q
CuK/+jH2Uk2J8QkriijhFj6xaIaPVq8IME3Pims2fZIv88ThVDwIyDgDtFYp21Dt
2Vupzz+eRKD6NqQHGepeqXMbMXJAEwPoz0PrGRVk3Qv9zY74UmzwnoX1u6cKlbfq
lzauVGy/aKzmpXevKmTja1oRPjPJbkrkiEtdfcXbAB6715jBBTcCFBSTSEJUVe1b
WdxlIE6QNQEn+uHdQn7ufJtru9KSeEXebtcU38iBGzM9BJUavwQOPR+fBhthVjn6
WZzsgj8P+7EEzAMUAiLvkElFBhB96Sf1E4Q9oFZ6akocSULQLaQtbfEo8+/uMMWd
xsXLgimOjuwoXPXsvSqx5tum9PfTt/IYIuCX6xV8kGx6+my0zvDLZbRUBkscqQ62
DZ6kVwJ8pms1Sab9wHem+y3L1mK0JF4plfFpJ6GTV6uV/m31nDaWj6Dti3MazeFL
HVLGE2G5XOFkYNf3dZsmJY7Xr0GElzZQ+5GrhaSAA5KUDn+RucqvZTcQ0nXexWX5
dCtP9lQhlu8eirw/4ialQvnOUYTp0MXwsXiZ1yUdTjEXSOONKF5Pi0cOXSOOXnLk
uWbActxwM4heR3X4fiI6//aLMvexfP242BEljoWvfNy7G7yGEfFq86dEapqdyZae
4DBKgLpsKPs0gJ42r7jpe3lN1le1GpV94n2NB1H0jFziGWqG6zZJ1hHjyVnKmXdw
6yXbRFRQQ6rkoCo+98KiTqrpdFD8YNKp3QSYqFQVcyqUfa8GbjyOCJs5mf5Q0n9P
tus/bfSf/S63JWhhg6/fHi6itceIkYKFBvPfOQHjRCU3N4WAGqO83agYg8hXPyzL
nx140qcVZK332O2JYM2dzQxT4i0Z7A2J2QzyUxN9ymSTBX/CDEaCZHHajBc0cX08
p2qStRyMHMX1SPH1t0UiON2ZjcgGxQRSYo80KWKe0S9Z6vaD8AcNyYlFzhyqmrD9
ZMkqaWtz/FK9uwIZWzYDuZZAxjutFwKKWSXR7rTZLT3wSV/BMUJmcLqUGYcHLm9J
ueWnlUbwknQL0cXz6uBHRmt/cgyFHBplEG2CP24mUThUE4z6e4SbJuc1/B9pOCB/
AKmUetyFzPdDdkixK7OzvPjM6zVJQAyXISHR60FdHMtHrUktqqctXqPkJ6w9fOhr
wq6QKnVNMyJa5zULQLQWRm2ionn0goRRBgVmhdoLH0ZSojDKI4HhjRMyNc8Jksew
4nM+VvmzlXF2H65FfAfwFI2Mw4LpSL2s17Tl7KaCQ8WgU6UuzH0p6BM/Vs3ckOLt
RxLL1G8SN1e2nhj8hWMAs2G95roa95woo/GXlhCkP7y1lzLIKkmExjZrHcytrAdz
oiUK5r5ctkBk0z1Jn4dGRw5lImIHgWN8oDwkl+USF5gENQCghOptX7uCG1mtkCE/
G3IrIeNP8MqxYImnuKXK8+bGYrKe0uQepkyHpqiTkoj/WiqzfL2j7WTcjls3NP+6
K7ndUrQC7fZ77JbjXL6Yb0fmv6sSrWrFdyNQeYkaGTfMyJRjCnOxzYfMUf1dZla6
w4IBDABx30944fGRIqzi4BmnxTHQZT2G6KXQMrY3nuUrs2KT594I11LJ8YxX+8qD
fe6Qog1Gk2mzpePgXr5m9g9VOhar49ZUC4jQFw4fZjJ+MuG2oM6t8iVqX3+GgpIf
bex4r3VYGFw1a8r70DaeMmjX5CqXsCExBOjvHEQRE5aPFINC+GWVjKxh9yFey270
j8+a1iv8kGHSFcrBeI/6PMheuzCarFMgAvWcTdT4TtvQBUD6RPu9nFXKKA0GC2W9
qyaiHvrtf2RgL9da5sVgXTSLCznPHYpNkyyO0b1F35PSNagBSjtjpsiTlX1JTqQW
Dq7g4iBYD4N9YcutGqmvED3S5yitw3Fe0NUD+0ysf7sTkBi1uKe3NAxfvSPwFeAl
znZAfIJJX5GX/KW1jdV4EMTcH2Moi6LuXM54m4FBenitPxyyLBtd2Vnzm151+Q8S
Ko95qQPLVtwC0armGalDvHMODrE9DTxhETrNUcZrHRsAGDwQUwxpxXhaDzGLn/DW
6QkOC0wLi4/2Sp6ZTh3cCTlyQOnCZAx8S3A63BFqEiwh5OLPsPZWpPNLYlUbMh5X
tw5/7B8UhGCkJ6jFNwH5mP+c0v6Ixysslu8nLv4zlIykCUXiR+6UjwHmLjaVG2F3
7Domwtf4q+YHn5OUeeM4hDI93k9LAiXs5amoqUPTTwHZB4wMaXEYCtTtjTQ9cwTd
AtfSpwpdMyp2K4nURAS+kZl5D+CGRyr6/vlKfYZlAVBgHSJtjLJwU5c8AKTerIob
/t78p9dE1gFu4rKIqxc/moWrYb/oom5GrrWi3s2COPuazyxErw+tpzPnWDiiSoXg
j3A43uUQiLViFqAFYZazHlQ+24FEnKkLoHdcQqbdtHaYZWILh6eJns3tLRwAvj4N
FjDDbnsiQOWNy/cksepN/oiwIhue9bglYJg44JBxoenk8v9jVN68PB/IUG8x+m5q
WcvfN+ikFbU3LgwHib3yEfxFxelQsu+D265NEZDf4JrydR74RHiOAO9hS4tBr4uc
h0da5MpYD1lPJlJJniTCm8t3MQyh9LUjjbTrfoWefZXdY4oAkWivo8vJ6wagiSt0
nUUe4CMswaPVuCrwInjpUsmDVVAuEQuIL8kx+URHDoI6SLqJJ+DyzL25BbUQGvss
miV4zn977F3YJvTxmI+Xjwi2yo1dBVZMzgI/fe5+d70EbLCnsl3/K3iTK4t23+jj
1N9GIB2wBj4iA9rSSK0/eQ2pUXGVfS29+RCczXPZeXhiUoEcnSWMiXG0gLJQbzta
F86ML2PCIhlQ7sN6v0RW+aDNcI2qhVOMdmZEZhNWZYdRHcEclraSzzN8yzBbI7Fz
NK33T626PWXnJGdwm7d/o7qgI8aFFrGR4nhM0yRl0I0yMV7+k6127rQO7jOIm8QN
4xYpt7SJbrTqg/smzN14/JYCtH7yoTa2lT8Q6SbRHOZazpQhZUY4Bf9Yb4pGbQcG
dmX5tUtJb2RoZVTP2L/ehLw/V3vxO/iJ8KvA9ynt1EmjWar9p0ZCeaHYqMVp1sa6
Lb0uSgsBrYsGqNDAmlNVzwBPnrsyU9veTzceimIrjhug/gWd8ujc+StAPER1NFNA
bn8qWda0kPwoav+o5g4t6mOHghgxRdEDMXVNATY7f5YI0v0lLyhJ5Yqq+1VxQh2u
ZygnPE6KAb1/N2nUvD+IUInuCI93fxZqvkcIceWaiOaqYS4sT5y7aUbAVbLoGPXX
zVaKnpenl8UVnx9kCyroA1LnPoi5aRejZ048EdKhNRquH1Hz+pla7osOJyzXSH4B
FZJenLzrHMAtuLClAS2tMcf6iZqd+j0ayJPMjjlreQSmtYzmAjZHr16CnlE7Is90
v+3nHp74MfsIcLouy3WBAiQtTOIzC/YL2I9ogc1SUBT90j5J/4GoLawbrI6v/47j
nBPIJwSayfZBEJXeJDJOd6GJvrU1iBlKNykOVS1ltw0/LM4OGbqYpR+062PsbdBf
PjK/nqusB2hlqWdavnRzUVJUIS8QtUk2a0NxRFxDd13+WCz7BPT8ba8iKEUjOxVE
5ahmdU+MZBrv/nLP8dr+U+gg4LoCZfWM13Wfc9vvZwNcHhGoFXQ/LY3qyNbxIQZw
Q9EaOr3IQf5J4XI0/8SESQtm3M2HeseM60K0QmQHeu+PW444JYT2C2PC4iKxDwEE
Ncf6i6E8Jja2wlEgr9+9d7dRSBjNGOE7mXZXQrHaXkX/WmIHIrWtIFI516UuRCTW
0zJF/RlbOQsv55uhTxyL9HEcPvp2dNeHrsfP9CjfEMxvEWTe/Ovq84t0MUv5Zrt5
dM22UtQjY4RF+r1vKTEAbzC/26HPbQ/nNB54tmooUdSPq8Fg88esxr2uqnihxr2n
KEQrc+Bpii8az4uxK7qLWaYY2LmuydF6Jjpxm3M2emrujaLU5L2LuHdvFlE/ncD7
WTraxmsqnFUv3RdtoqLU3qTuvulPlS9meZsbSFP++NEqWrEOp0PTpKNinbJr1F7e
d6lDwZOUjv3ZXqgTDKY79SE/73IGQW4u9Tm3hjHkzWOQSZ7Cx6g2xZOsCUYJmOI7
FcRT6XxzyASC84915sGrSANS0OD0R+otzNBIdA8+MCfMXlcjJJhccbtqU/znEgAe
h2YshGD/SdcSnbFNcxoEzzvYeyhzm0pVPUew3WO68iqX8fGmaz8aRUKlRNqNLc/p
qJO/n84PzOuOlvKWsuEY8bqY0xehP/zftM5g5F1Y4KtUI8tPqjth4y9FJnQydSWX
X9TfS4MT+l5cA4eicu3l8Vdpbty6pNKSkUr+FQuuERLXY1k4SvatYMFT+451MjKU
tvh/Y6CTe9oG+DW9YUqiyPYzXLwn/QpPYlJabesK4uKB01IxCT6jf4ZjRn+9FH3p
xVCw6HpdpvIwizwE4wf71Rhs2BZwh/MUFVkmfJvHucpzSwXzF+N/lEGUUZ/2zBHN
2ZfvZ2IY1hPrWJ69GXKlQrefqby7vZc8wGA46100lz5WWkC5/q6V/d1czr9UyLIF
uCgxgQV5C7bBqEY8pANli1AvyKMh0BrtGEhxc8z6lSlKZOzRqH5Tb8BgMfZXaNQX
o+RrunO2jwDsY/JkAdKK9H9Wn2oXvFdHryFyWOE1p32bjkbguDXR+5UDsXuhFemt
WkjsDZKHP+z4UnSUzjRDs1YPwAfr1riWgVERGuoHevPq/rTfE4FY2UryYuc8aknh
QMEW2IN/jv0peIVtqmxomnJ0TVXfkfVcrjIrUWxJ+9M2pFLCepMzwU3va5X/I1oz
NoRRj6m69n5UHLsNbDkEM3F/5UvUv7CU/aGce9nYYsYg8mRA6J+fj6VJcuggm880
iQDUUJucgLJ63srl+tmt3Kiy/mm6IKY8uhCgC8f+ojzBQsYZ8EeMWCGmIPqcP2Jn
1iQq6ocTlLud1fsmf4fRXg5dar0H2UJ8zipJiejf7lxEl3zjQJpjZjsu4BIAtkq8
b5Ph8ThZ4iYWnz3v02IgSC2tuXGqgPHscqtiCx7wVTG6MhB47C49mPhNhEVBGM2u
AkYQfH9DANjnOTME/ecFqIyluidMHBoK+sGICZyuxFefWAuiH756p+C3Sq+OTQqD
We7ek6WeA5h4ByoJd7s81wS5EonBR/ZsEAS1uf9AmEEOopYVzKCoJe22LraNvYb5
PKw2sr/kNORgvdcFfWUoM/GsmncQrjVUyACP4AjBmarB+bEc7C3TzAb2HsHF/6lq
JV9BPgicUYmQ2EMAuSgrDjd1tV0tRtHazTZzT1bsLj2huuliaZtY5jQwYGzJ6dYa
2yavAJpuggyM67yHVDKAcu0rrfDZarl8YcyS2tyDLVloOgS0GVya2JMswTM0G8/I
49hd0amwxX5nClC85MPscEbbdhhGOkptm4tUSZTBJAAR/6xjC5GxJuM3OJ1+IHgA
qMaCe0UIK0LtHu7eF6Kub4I5sDJ8btKal3JSrJeu9VIEjpIwq6b7kcu4YtOcudQ8
zQ7gKCFoHsDXny2jnRQ1LRr/KYHh+YJa2UvQEwvLUsAL2tf3QW0fzZX7kM7TXjVN
Ve3TJxDs0iouJZvQwcbwvvFmJeAFE8QtiyjKAkmMESzJfsMQamgHg0Ik8x89+T72
B6N4ZMjYGXKn5noFzxw7qqDaYTEiXeEYNZjHLGSA2gKVBCg2xiFoU3eS15LjDVk9
D83qIwYI/1l94u7XVpqPtEDRKFGpQ6MB7M/PBSxftChVuHGX5bIVh6JHOxUzTFDl
EELifiEhwkhavSpioY/spNPed2xi9jJpO74x8CDPDNtRxgJW27CELtQuRkSfV4Vj
sa+R2Wf/WcfIVlCXNrHh/XtN9p0T5jw+0g0OWn+dwytH3P/r0oloL+sH1b+9ZyqV
38caL0JiFoKF6PEEhqCVfqsii1UvPpcp7+c99kgIuFjeUDj70OG2KF0YQcPS51Ay
Kd5RFcJureQyvi+1a227M4MKwniFOHfHUZ5oPLNxdkiS8D21c2WGc7WSWjCz26xX
ROMfqjnikz9vlNulfLIVFy24Xlk+ZPbGA6Xp/Me2IrxmN5npoaLCYoJ0R/RpvjMI
Euj0K7eD6s/zVSclcUobL6NRpBkMirfqoCinkNjEpo/aHG/8xePfuLeRTfnngswh
KWohWHKvI1q0GSeE2HBSLQrwTmjEEPDBffeOwmp6F/64qDoXh9NE2kJLbU7tXR9Y
y6AoWOdyxr9uuhk1IYJ5DPMy8qUacmxwb4thFjxMAa3CTMQE/NtReSIeQVg2pmV2
fZWNcVCH5/EVc3xsFolUJ5xssxeat2Ggy+S+UsbQQuWjkHZbiVO+Js2nE8zREBnb
XTPYQGTy9qnH1Bjb1OuWfTRBBwE6z5Sks8ILWWQRQNT1Mc9ni33MWeq6ECG5ANge
ieUzNqJE+RCGyW/5eEEsCzMOvHWtVOPzlfsDAq9m7VoL0io0+E+WquDBLoq++UwQ
f3nsW/Ye1l5Wlz7R3QbVn35EKM9y0+kJbLAis1gFVWvZim409PNA6rvYBTFCRxLB
NZQyaZkvmPtb1wTKtygBHDak6G8/RGpqvYYXQQUN8VUHMxbTsQMcTxsDdv+5tyMC
6K0ZsltU7ynNVIBst/jFgX+Cyda65eoGu9UvF8jmFvnHLbH8LxFmyEPbWwdbdsj+
YHsKACbDMIEAhgtSoMqNTt4uoRJzxFYy6RvK+jMJCJOsqp5/viaZLsDvK+McLd+X
4pRlnn+ttfSTy/6dW/dYKgVim4NhQIIggj0R88Bf3gz6Xq2yYsHDfEnaQxO6OCjk
q57Ft96jOm8H/gc9rdAObS/4q0a3uJ/9TxPqjKBdxK29XqhfI7wHFkTR21bM6CXO
lxCkoywmYCGYGMjqTJVWhg4ETAcd2AiOQSXmdq3XYb1Lo9tBQujXuXI0Smos3Wfh
r3xZRofiOwvS0t/r3BYDlRVVZZS99Z8Kks2w9MOgTMGtYRzW2U0UoXw2fvUluixS
UNJicMIfs/DqIXKE9/8VmT78m7DPhF/zHv/kgyK9mZDdTyMQKZ+TJbZpqHbKJZge
jBg271MQtuRLBn04h9OpjXG7ESCa+L+P+YtwBWdHD8wr3hlWEG5JsAybDCqlxY0t
ra0F2iNPJbVovpq43oNsjuymk2WqVp8KJ1QXkPLgXBuHsTWVGpwYartPXKcxBLTo
2gk608xHxfTn+lTM8LhJIiBt+up3gM4nU3VFCkT3D6NSzIZrJJxj1v8z6REajUdG
qebP1kcLJKMvJEFm52HnVOUktkBYtktYLnmxR3J4O4ACZgFOGm19LEepC1gSa9mw
GjQ8G7UB1yoI5ryicrH33w9yB4jgde22fNdYNdwpnFNW4UDc1bMxPdbvitKqvMrt
kuePheYIY4TdW2B4MsC53kjG3s31TTusMZd39Q/iaUXUM12vXYgPhwgS1wIyeuxq
FlSUAxCm2Z1N2Xm0qTfZPviGBA/MSFBoGGeRYHBB5Gw+fPE3V6IFzTILtzy3alXe
NAyrAWyxhZr/X9qltJYyruUkoxQ7pZ/m+xSbXldpuDIj9o8haa8DRyK5a7ogc6Pi
kP0TtDJ3K04DfGvuk0jurY+YaUfCUqsCKrwdl9MsInvIA23JNUskImcpWuG2PYDM
b3Q11kjs5O6VXoyrrtLWqM9Ewgv0GtnRnT8njgyG6CPWGlgSRhBHI44eyhAed9bl
UngLXW27Nir5qGmrVkoTYCdmfrQotAr+b0QMRiVZfxxdC+ZsSW+0Tw0IBmnNipe8
NOf/fRoOWgUbVDFTgOSnwPwi/KDYgwpPN5b5eLwkTDRNwEcf/h1tzL8qC4V1Pa0c
AwP5yMJtpNagkZZin/WcEGLJt5xNH5gtlZdQmg2+0tYmYfURy/Pu7RzwL3KiP4oh
5wbxUMQ5cdWiJRyWLHuR8ztpvsj7PQs74EeH/396R9/0uuPQDZ+lFBGUzNDWP24w
LwZixSYhSmIV3ywN2Wrf2wYotfrGXOh2Vfwnc9Mepzxyia4tBjLvBCEr/7y/GNQ/
bwXtUAX2DE6GOk8n6TmyLptIBnNt+CrVu8hXJktekRNQT81FGYGSN9+1U/EqOQjr
zptWIJqwEf5dmXUccjTH3LX3iOOwwNbJiPTQF7JdFHVRFwd78wT25bzWYE/a8rUb
cH+8q88y9fjSjeXSYBK65CkFqLLzkHH+ZVq2sockx1OmdWPZl6DOzzImXVOLditT
mGPY9dw/zZ1B/OaYhN+IK8ZdWCrT1go8zhKFulziVvV9rLa+OhbDv8ASkvcYHniw
J6pIUF03yNAlNuuU2oCcNbmOQfF+sHqMqFsUGGGmTLv9XqkrjFQZDaLpiA404zAv
h2FUoDbkmCUA/M1M+1uRrc8Ad1nm2ZGp+lin4QVrpYWTX6arKsk6gTGaoWbRnRo9
yGTtrOs1xnjjiO5J8HqXhTXbUF4BR62qJao/SoLoK4Bscfq84boUyFvIJ36zTNud
lU1DKJtGBzXl1PjW2GOZBjy8S/bXAXtT2bm1zGrrFm+ZbZuNJ1Bg4NW4LRJv2246
mkLGTpXVjM8r+7CNcV6y9v99tUa6S8NY4+JSEhc21jAmA5O1RpFJzPNLmcCThBHv
me0B2cD8Oq0Fzq3mUoyvKVgI26Et/knuSECvMP7CuvVVL7HyIXICJDso20M1I/u5
WobbLjyn7+3Kf6YhM9pfYDVVqN8wP3xX4TaYAONppphuIghDoOOfQ/6Qo9wYt3rw
Wt1duv4dSBAxvl/xuvirLAzXyr2vcgw3z+3Daf6iemU/MgQyLPeSfnA7/D+DsXpS
qYtK3d1kbzX9FiT5otkt0JwVglYxyTnYjyKylBPeLmYHiq4zbZHafJ4zKdrssoBi
XyKskOjhxaiGJSmoqsuRuh3b5XGknDAS54mMDIunQhzlOxo5YfDETPydJcxfn6om
6LaVxJuo0cUmEj20Cs6eN7wrBQo+Oxore0ViuCpAWHvr33AdwlijyOS7wc9xv+Nf
8c5M+7vexP1STLoI5d5OW86Y0krirFlN/eT8q3Qd0jeIyWOaySym94Erkbf4Nw0G
NeoGEv7n0Puw5aXTpbb14fuQhLiQ+HjVXXsQENW1bJS/U9ZhLazMxFdgVIbxxITY
/9aNjCKdcRc3TNqQdXvij3XVey77P8cCkoD2fo1tSTvJgGWToj4hixcPUucNAO9E
djJPpoaxWl58+OvIcmqd97jezJIOy2EPjkROhS+PL6ImCiWah8HkIFhL6bNxkC+o
7HQlGMtFeNc9K44hHPMWVPHv/pDTvjmN2ZlpzFBLbzZE5+23y9be3J7n1qmFkEn5
KKAnqH4oHNMJFhA8MvX6iRBWFsqnOsHxg14Go4+KuqEjD9aQpxs3rCuiZ6j+JIMC
QbM9lx42qc2v8K/k1hN3nhcxWwe9ONy9Aa5Qg5NmcsM1eHiRdI1WnZ/vpEmp4VXv
0SRBIGpLyaXcWeoXSnl43E5cvjDpo7WtNTac2reowY7OFdYi1YSM8BsWmuRGbIw+
PbzobQrsi9viJsN7HVPtRv6LlOFcrpdYZl/5/BzP+jf+2Yqjf5itHxvnyE82v7sr
JS1YTuSJ5/vEmFcp1d7g6iZHN/rD2Cu4gmaRW/2x62DW9e2W96eJ/z2UZKyeJ40C
eOF4AKmPSgG8JcFRvfVsx2tcwcvT+mcfLNse8TFL8AdPBVzkMFvPltO7rL3kK9St
FunXzhO5ZcN1QwLRP9OEfoOxM9a1Jh/YOphAc1GibKOYjHz1U8dWUbKtmFk+RjZo
iqU8lXxTFEl4XJdi09T7xS2FoYASWC+Nqo2614rUiiBNezDJRk0azkWaH3TmuI5C
jEAXZbtmi0+gtkbN/LpwaD0L4oedjNLadt9obeL8N3SW+tD5drCNuEADBFMEFUAh
7D4OdHYK4H+cSzHOtVmFX2bTtt1AhUz1hnx1C5JKav/QLNLMb5HTmIpNvSHdc5i/
O8XJUfi51rcLJcXH3WLi8T15OB7Qe15/C+ZrgoH5+k8PKwln/UZY6nXbuZS8C9Ry
oVPu88mRYL2Rc09nwG420B0snpawWmVKxzrPkWM033wY9helWsuG4pDUL9n0Y7EE
ubf5L/d/rHAGX7dTX+RreXNM+OA2vyfSNi42YCdHElQmS7LoIrwN3EodrK3Z/HH3
BIzhH52NkkFKx4MSdTUfN0Uaf6wocLwDvyL8hBTjpEf95ufp3UbAJv/s1QCol3hT
G2ZqcsWLbFhTSshZCtJqbhK56SfrlYN03B/EwHDpUnaeN40vf5rQ0ePhHs4j5Jrh
AQFjGTlW0dwOxjo9FQHRYnoXE81wrnBsEOXOi9JpTZkMLnyNfydrZToDbDJdV0RD
qjHTdJYolyGKpb9vp07Md7w7FB3f9Y2uuLm2ZU5soIK5LH13PJf16ssUwqeYpLBT
zvNf3352bv393wqy+b2OmKh00WhCN517Fz8wLsmgJi/Lu4Q3+LsTqjnVPKFmB/Gi
1lmg5XfsXJKNt+CR5AYOgwIP2IsOWcqe4IADLE0H5LR4+6CbQXha4C6YfkOC87nc
cvls3kG4pdeVlvMQSYFCEilb6j1x++ZPSgosQAbW+qY7vVb8sCx7Y+0oHusZlp0n
fgB0qJfEZDUJYNeqRQy2cTSLgK/hPPKctC2aSJXB+5hkRLKwva139DGm6bBJgxOG
EEib/dXvrVF5M/nT46F8+PeYJu4FB6qwaGya6Twu9TnDwD3fCTLIn7OilaJ5x5MS
upBzL7S+CxfB/IjsnqBsGuuLKJjGtCWoDBKNQ4xeFqv/JzgJn9mJnumm9QZ3S36X
ZGXzXX3PxsflH7RoQ4WaWSj4gXKmujlEhJ6CEUZJixNGVOzXJrIsnkFEBkC+jhBb
O3yjp7Xqz8RTCpxQ84t2tMszfE1MsT350hXn0T2iQLMjr0RjknnDV3Ofl0OSoGEa
ovWeEYwzDt3huUZXxLSxi9VnLOKT5pVGfxpKhqEIcXoYr/HptGaGjq951HqsZzwY
1cEYglFw4B6d4VRlM7LQYNeBBoObE0UuqmCe/wOAZwJilGXva13Sf4dHiqk0gM7q
kp9WzxSlD+7eK21z61AQMZsz7nFlK6ZopYeLpJiuqGDRlS4j0OOfHM+FiM5lfxM+
pLh9CkMZAOaXLyFpWYhR54kJnPvyPWYQE6D1PKAizX/yosDa+0RuOnfFJCx7XEzx
TqVaiEHp9aipthQvrn0+RjZBXRMaF6tVtwncdNyo0G7rSRSG78AA1ZaQDlpujsNM
fqCrfOyJVQFzqsZQL87UcG7RCcJpltFtIDxs/8Zi4s2RPWNwWevE0xt3BWIGT/V1
/sYHhgNYj30uUkHMm2bFV6gWeTSgRA7mdnDgLdlZiVO3cl0JrkRIp2FOcU7c/uP/
Y5Zru1LyjXb+z+/4kz5uuGG+gBHS8ULRBZ8d/JwVZA1Ggd2QqMX2+Sm+Q/YLR2ma
GlYH1Lw3EV3JkuZJSOLYXd6msuekcXEa5CWAAXt5FaIVG+uTlcxfIkSBXK7EqbZy
mwujDzlKKwRR7x3MzTiHoLwPsjEMHoVi7apxROKbTEnap1UMOPetNaKb+jpRudOy
DKrVx6g5WKMADHzIWPAjblvidiW/J4/HTHyxL3YNpEKyJGFioXNCV+c92GHwnM0j
3IXvGDblnSXo1sjruWbAyEHXQrp4Em6Ni4sL2w1M+uaGjfJEcaZpoSkzlFV3+U9r
ftIGVy8/fI+cDHuCXDoE8oZjOiqbfGdyVbMDkEPLQDCkeSovMrnwIB+qcEbr4ol4
kBthoRAkYTPMGkzWL3HAZSwmX6U3jRF2JyIfJ9bh0bv0TPudFg4li3iCJMKlF48c
0uFwRcAhrsxcdvFpfNjxBeEYs80fYyZt7IWycnzCj63L5TebqGEVO8BGV+9iFwAo
9BUlvZhHc44QOPehBgyMmYS/DQFTApxXgae2uq07930kWwQnpNiGqk88rus73n9/
lQM0qUZf+nAYdU6bcaXhcN/MtP5z/3jL7IWkqkrDwhz3JKJjIqhZx7UIssuxCKD8
kXw8auEngKZZi1/R2VEDlaQe2yY9XIB8hifrG5l6xuvigW310ZU4O5VNyk/ONg2u
gompNqLJQfpn6Vguzt6kx6nRmW4RARLsvMGjX1qoM1XQGZ5CB1vhxhih6QMc1QjD
YkzH5BMK2NrQK1ujRx2yyzN2xelPwB98WdtlYALqOLTYYg7NzPu6HPVCDEYnHkWH
TK4N6OzbD0NBz4WdG2q5Ao+n+TNEhVw7qGRfrrIRHjErP51V5b1LIhzZ9X7WEpOo
vlaSx6cwoZEyw1tBY0VYafA9XBExPXLw6IElCr8D4AgPLGlqAbGXcQ3BVBdMsbBM
qNqKPwQLApzcirKH3Rl8rE0hzMaacHpRdiHOe/1n71qjs9Bdxa8EOHWlUlxLs8rG
SeFwOF7/VnzKozCHiMP7UnYJHGIPty9QB62J4ZpBsS2i1/urFWB2W+1oW/uuRQEv
iOaVBG64snPxZUCNeFEBvaEPXR/2/kbm4za2EJeAd+nWf3jda9Ofr35n/prrVgqF
9n2SijN7kwH+7q7nd0Yg7+4apyIU0+jATbwdSoYP+7PNPJMvQUW2cgUCxJnmAZjW
HkpKnNn9rG6pcx3X8CeAuHP+ADD6E0TIQC8OtMkw0anni24K7t9nFJoYKUmNEAPA
kEkHnBaS6RCeFHon+l++vRwhVxg+XX9BzngmIHD0inxhes4+3dg7+6A9SlSOws+3
cr/c1tv7LChtw+hc13ksCIt4c1htjnI6aJxx240OVnIHTYRQfYn9O9FtpBlc1QDB
UUrfgp9Q5S4Qv9KWERsF/cbvH57q03E8VvA41u+80o9ys60bKrZusuf8JiOh39Yc
DOMzrhT465dG9/regDTM7wCK/J5ureTPWDav+QuxOnpbvDAsUEdt5SjgGr8csXcL
d6dn77KKrRpayZDbClnwSXQMRx/N/+3MULOG+DKCtY9/Cr/5rOHRhdymsiA9HGnx
uaNWeF0rHxOHLxLW2o0ReLHXjrZSDecfbfupee6TlDQjitPTHBn2E5+VGpJ5GuLh
tVPZQGevD+AhaCvbqcIxGL6mUnz9GkoI2oNH9DDNbb8W7yzDrM9BUTASVN49nus1
RrxFxcLOZycKcDM5wCvFmFSK2GwGxoxWz3zfC/oY40FArrusKExxYiJrrhWoNVs5
gSAB5KS+Bg4TdBD2n56a5rxTnsFMqAZIzgPqLT6viP9UUf14HWizNrmqSY9SMEYP
vvE96LHFoXxvmF2epKk9KFXcXNv/LViRkEc3vG8r5UA/bsShmHKwAj1jtOPCKPe4
Ou4LOscN190jzjWVuAebEXOOmWA8IYd1AIwcjTZErliTPCPcjmuv3iiSDpx/7kyn
X4Cypr1UPRnOL9+0CfTFj8Kku9Plfj/00Syk7sib0mCKq8+vWlyz4c6fU2+UPyv7
JJ7Paldkfq0AEufT9VRIZCOWHwywe9fgwxuJVGxmfkuHWsFu/+0WMecyuO2GXmF4
3eArU694/m7wYNIDmCLnCFc2yvxxlUNVGCrpAerSgRX7BR8q6TjsfyM/wu+mFtDs
FjIE0Q885oHeiHF7VIuCONAZgtomVRMbEFXdtP4zUhq2q5x/vqFHoR67XzM/Duc5
CPBbVGhjfBChuqu8xvsR2v7r0yhc3MmTj3ejbVDMq11duh4JuQu/A6yx2xZg+X9w
INAIbi0cvVYokPKwCguFPEu2NZKePyj0b1gCSWyI4GFVzjUnAjb2o2KVtykWRHru
iLre9PObcpxEd0v6l3kI9thqrzFhXIkycu4QhmBDZyDvUna2Hkgo3nsG/xsDM/9D
qge8LgoNn5lGZqETnmFz9WGlEkSbpfuMEUY64BfL2ySvdq93xfUZUF6DJ9lOBsCQ
aNIa2WkCw3XG3zvRPx5zllRiP2cUVLra7yDP508aQ7/NpALY3n3kkAL8LB8zrJ6z
99EIl/po2T4411NtmCm4q0y6di08egxSCqRAPjHhFyN7zO/+u36nH4ZpPFsyUwrA
uT1ZV+3qJGVRB8WqnAPYr/EhO93UDYWntNGBbFCsdXvOEUwEDcxaXeLEPRgtvMEW
EhrYsXNTF5p9esrgac5dBPMC6ORIa0i6vKieRegc9N6TwJHkzZK2wt7vbvPM+Jqg
mhXuoCIZdkfnlHrf6E+NNwt0ziMGGqua7uAIBM8nkPUdF17GEXnNapMwiHKRAUHB
yRxTqv00I7NHRbQ1YK7dNvs0ncNJk7Ns2Uf4SuPR1pgODkzINiYeAXahcHGwbiGR
cfILmvqSqiG8y3KE/PfPa8XoQSRbNeD+1Xz/FyFBlxcQmF09mQ9gAc14hrpDu9qH
q3GQQT3JBnT+pzSON3tRSbj9Ngeu8JVeAPSmb6iA3Zx6kll8sCh6+oxkEUOxz2+Y
N8ikJ8cru/8EecRHkqXsFTG6qmp45jF3oOPoA+ITjLDucYVwbU53hLeFNW99zroN
oKSF7VlseG5XV3Ko1yDi6N2oB3tagJShX1gwLyNPXEWJdP73ycWzLn/nNyYxtA/2
k/k9j4Gj4d1xjyXFAs359HL1DumO2MaKNRPW2l52rlpTJg7yWi1aQd4qoxcF4Bh1
UTRmdhyneWerxdCqKTN6mdGrNBmcpsHJ/LQsgWnueYJ94IoSlBDhwsDpcQsAFMDB
OfqFIJnzAvZoTDIk0+Nj8K8KTI7dHxP2TF5lfMsmomUPFL5Ltm8vO75PY0Jvpc43
zMNOxpRA9musEQP5y9qdvLlVd6r4jmitHGCzYbNV8gNMZMD+A4Hdt5jRKed8RSDs
+sQ5d1s+H6KmlMB3HbMxQMRv1sWi2t7EDl46bX8gPIbJhxNQJMPkGyjA4tLRu/vc
L6JSLjS9le7FtI1PR5z2GcIIu0kdXuul/q2CQ3LVDXh6x9L1Q7l64MkORqhJjF8u
KPwWBcWEYNenWr7RFYZvhFu6KJECDEHx/Al5rpnzTgcFa7MF3S9SOCYPd2GI9Emw
mbdVMkuXHvco2tbniu446Cd5QQeyCLVokQvzulLoTyP0Ig5QVmxUWhvzifuyESJn
GpVH97woM+sCR9TcnvT+Y0UOB5SnVrGPKatw4KkNmvzwdhYLKNSW6Bw2RMv4cwfF
cfyDgYrHza1w0EypLTHr2wdC+Z0NOWHJirhphqjqN7y+ZajILwkpvFXOTNWvhBup
eIkG0P1sgXaGLHpFBTJ+66BM5cqfgAnfsqDFXCdBjBHaCqNlJEn6QPsj5ni0drs2
jvsFEMTzY9pFXsZ2dEALYApCL3YNaixwy2Act35RC+4XYHY1khEd0BpOw1L9sxtc
Uh2Ag1nenFyn9vOkimdYtPJXBwGQ3NuLw3L97WTdcbYd07byo/KnYcNi3vm0k8Z0
wmiid2In0R/wTBPg9wAf+94kcxHw+BXqOIyh2VQRODtZ96YFwI2veKcouTvUJmou
fUmdE6ROKOBkRV0fwBXL2vsEKozk6h8Dy7Pn8ZJqtqQHhNZXE95dhtw8HBqdPqS0
dhasJ+3cOrIOJBJTUNtqu/xAE1Hu4SwIzsFd8xpqrY3eKqM4DZ9jLXTiiGz05guL
yZCWfFwMmb8Redq63/Ew/DAJ0XualQuSsstCyE73+gh+PbBG1FMkZFSQdkqsW8UG
eJkpjyTdwUSjSiKJcLePiOwYL/iPP1W1q5Ai05bvYfqpUUdzi393h5ZJG0xqyrN6
K49kSmzFOd84c7U4k+BfcqqYQ7Yz2w7+sH5xSy9CvcD9QHunL8yGMsnrPxSpkMoK
fivAH6rmTEPRRge82DXWoRC/1s5Y3Dvdct2TBxSXqPH5qiK2X4vl6f7Up8xZifIG
mwDC1erYTKNmeeCgJ+a13fx0EjxcZateVUF35KVfo2KOoUHEhB0YtH7tj8dTjLwh
LpLW2Z9VOEwP9cnGSHP3mOVU8Wa4EtKlelF6wx5RaiO9wsYjPbYfny2WGz3FBpH5
a1YKhp/x2HYsgjpVL+VKf2adBcXUF0m/L2sf7iANYtmFpS4qe53t0piYo3fWEJBw
2cCGfeAlvLjAbDuZEgPdGyqIjCMh+t5483At4qYq9W0DCzOds20PGuUqHx2icj7n
IqIs5lL1C0cBneoxZXo09Df8KnPrpeVmjHJMar88JJJRTX8eMROF56UkPtlIYlSR
S1pEEZeWRTyxStaZKT7HVJil7ouKBdRU6zJy9tn7yLRm87qW6TPLuIfLGTyiwfgu
NDYH9mMLNpNDJkySjSXzwuFpBKOAEzdDLnGm+w2a1ZPIwWNw2nv3sUGYxlKwDeCB
qa/mXB2XIwwEB0XA8Lgj+mnNpPrCOaiLtOJPpUgXqbp379++4U8RFVMggQv/YtbG
E0br73A0OdlH7z3YG6ZBWp7w5P9SAvpEx03ONwGhtwa7/MoFrZNDLLU1oCAMXAGA
pfdWUR62qYvjshInZ0S43HohoDiPJ2F6IvYnZTa3rH73BuJQh41gpKdijiFcS5n3
ZSVdtIDUdD7wM93NcaSZg5USDHokqMIGcdp9Jx1Wv5H6552fHB9dZDh2fHIPkVNu
u0mm5DKU1beplKmqrPm2ypUiOHSuZxPUrzxGZ1yqUBwD0JHuvKtb3Icjp2TI7Ul2
TXkMZ57Gw+JdoYRQ3x2To9iAFo4ZC3kPU6ndNS3r0gJRAK7aKCV2n13U2tBad01/
djITH5snKNbpVoshUEZ7RL8NA4RXrgRz9zHo+Ve4q2P0Zf6pNMG+mj11pgMcYS6y
cqIEGSiul5TpZq/sU1p3GQ5YIGv/4uaGV/VDstY3TQx9GKdxekSYDYzY/1xyOE5Y
PFIIvALeaVP1udk3r21tLrSUdeJCagp+spJQUpJpI/Z8LXAuugtvhbIAM/5d/U0q
mOM/XT0gtxntbVadFcEDBHw9aYBU3Sp2Wt5gwxFl69GYu2/g6T6UoYYxIFa0F1HH
lih9hDuhV1acjnlGJcjK8Le+PPfv/TFbbcZL68G0i6FnKVNurjjSIefal4GftQJ4
hkgJlYcQPtxy6sNIyf9BjEvhnUHpxRA3kYUPW5WUnENMWNxfMk+yY1+ZxU/pSWZJ
JLS/vzxxfPHU2svpm4CO4BXdP1e31cI3wbuKqff0UjO7UakcR8mR3KDym1S1+vkl
hK9wxVwAMvFxCm15oJfLMyN1xqagwnWI/TgY+hnZ4qMqoKdjj21MgbhDh1IClrTE
8Rx45YeoaWswlSu4SkcEgbGU+PiingmhtXaJHJ7BtrtXfowHsxwAaPSX2iG2oOMT
69jAOHGkpYdFTF15nPaegOC7DXc2Wv8qc72epBSdhSNicR/Qay5AVyyfOzDlISQd
SLPmlBaYy+Ree+6+h9TqlpuJONpJR7Xajn2lo5/arFgxrKqw1ok1e2BD0Vd+7fBs
/kKvKXrlH4ape5CMT7orMkSO7jlLOikWvIQTeWngNCOV83sC3/fEIkg5s4uCpD8a
fIek+3fw2YXGV8SCGk37FQP+ugAStci9BB6rproltCtFm0J9FurLb36XGzCXNRES
AHzopo9bAud0kh6BFw/K9oeRk50HcDseA5aP4P8dLR33HJFgXhQpjZlJvdaDnUXy
fZTjlIqMjc8YEoiIZaknEiQe56zXwaUKXHU4OF4ix0kVcn9LJthUJTTl7QBWZ/hg
FboUds+e065ysetN6FrE9ptTJujK2aaWaPJ4D/MFRHHtuXma4/9NgsgDpLaSpP2Z
rlzNvYfTzd38yEtP5gUFbIKjgc5Qhx4TTeRymjY2PhpJqI1pQf0svpx52JVJXOIT
xBEdA+BD94PeMx7ruajZhz3BtMvftGo2JNOEqAwMLS4bUel1gT7HU2u1wXahZ/e+
CjG920epzMtZnYnAjwIWJxzo7OiG/rJa2EMGxMo0dT1jw+Dk0UQ7fs7OUm1SmHE1
I0bktGmnYUybV7bTWXmLdZY3Cvnhp60IbbhPJBMjp/A20ngbEGdkPD30SUa5B5c2
l0wDGjgsa4Tu3wklS/oId8LIYezSAhj3lcnj0JTDMJdK1axMAR8gXRyUtnC5p8rc
IVqYeIDaTTVDDXGzljyAANrX98iV6jcfat3XxXa6l2waGlWon32XkWfLY++wC5rH
lKzNGX3Gi2Vw++HTW2jLqHHAiQnF6zGj9VM0JugwllnYz3kLazY2iHbVlkp86WU3
MMmRlDRNgsqsqQ26iLNjul7FONyUw73wlabGWGxH3DoS9kVvgNgjIiEcCBn9BpUE
HDE25ZZWaXfX+ZqTnlVEEvRs/Qvun/TKLV36m1YKE8ZsmeRiOc9ESXUJeTUBRD6Y
pYfv4yZQr9egw9P0bVeEvuBYaPFpJV6bilGFvNCIItAMuVureTG2ZejFNCn04Z3w
Ge5AuN7jgoiLY/scGzV8YQJLMiqtbS/FRfrIub86JIyoQBcthxY2gAoGYhuuEVeS
p/I52gDUjNJSWTiKQEtQMulIFDEcTd18HfnW23DS5uLY8ii9L+Y2hYmGKoFoU0yo
RMKG7zpd9/+d+NK8egT6rFJGsr/Aye4GDFmW3vHxFypvNuSyE7O6qbUdDRvMh86J
sWLuNaYMgyUwCdTMWT+LXCt3lFri0REnhK00iI5taDcsNEdEPfPRP1ycdd/Cnqc/
D/bQsd25JRf3DBxWSsDNAhJeqQ8FIuFJU5JedcRAppI4eIbL0/NWtVxgn/pcoa//
RkENnTGgKOvy0LWu4PXoW4HvjkPYUXZsQUo7ZbcOh9joGPQ2+BRMf3vrgLlFBYON
8z8P11NaG3m8utxND0LL+ZYr+HkGbT1v7CkpJIzJ7ORhBQ3Pydvyw+mApgRgSIH7
kOFmRcZEBGfQHRjntHNw8NEbh8q4L91M2Lk7dy/R7pMVNQPraxRH9gOZ4KBPMhGJ
N5ToXRMxoFKisrWra9u6H8CIBH18IhyKAHpgwlBVzUFky6nfpmOan2APIeMALVZQ
/YXI8xsGn0GVwiVMmEg8PPyktWN5qRyTGUyUJYaSOfFWIq8Y807xpM8SSeD7oRDS
aydF5bqQ6MZFRNQKOtf79Csny5YPQa/xXu7ZtRU15jfjwVpfwV+cOaeIXxOnSkLg
QcU+9kdXEte+DqgX4DUyRX8JauAqAvB/LXc6Ibc1NHkMi06Qx+1Y44BZ9QcaXKpN
1bizEmJLzo7uWeFpuypoz7m+c+p9um3hbti5ezVcAqeXPzrp4fedNOUAZp0SuGF8
yARCFQs400IDO2jg/69Lo1sSqd614A0HXc/NP125rE3qbeOQ80/5KIcrBKHdlG/j
FZuy++9DrOC9Pfk810pd8fX1hwYIg8+eF2Z9dyS/JckXgrECj8jvg9RNFhpFMttR
eMJFkX9w4qpWEhMCKg62OBfoODWzi79FWGfE22xxNu3NbD/Ztgs7h00Tiub9o3Yu
0p87g8Wjh/FwWdFEADVDK5CtC3L4N8c0bPdQJcQ+UIFEk0G3Ss67Sy+oL/H+c20N
1oEWo2Q7D6dYhrikHJ5TIRaqaCic45ZSQTrPGg8sVcQex0VYHIFkRr74dzhwmXNd
iEA+GWAlRgvmo0zjLaUUpizK1Z4cBkAdI2ZvTfG2cQtdIxMKrbmcG0NrDQyfvUn5
kvb5dbc3c2IKZ1c+am1paT7O+j+y4fZ+kYbNJJ9/OQfi+Uq9dah1dKA+0+XORp1A
et3ptni4PM1/gG+CDHuSmU0FrRaZL30lgBiPBWlHNY4fuSuaRohKdG11hkcAd8bO
o0SgcneZ2rGkulLbl7VCnUsqFH/kllNmr8C2FzDMbEogGNlkw3QNu1B40kzPJmuX
RK/BZA8XF9D/uYitJkfTJeH5+EOxKWRb4mWnUoG4j7ahyEnr8AxpMZlWC86lxKWN
RdcqJc+dtCT9duQSq9hQFxW29WwaQaFcyCWmeDfPDo8o+s7L5ja4xJgxewDMdS6F
twQZIGSXdMz833cqfY5eKnO/CBioyhsuSp2z+1GGDgGK+S/hpe5eSLQphpPVKocg
5UVuVl5uScapJe3S05Iz5lVNq4iEfdZXWCZBZbMRHMCAqkzi7I761G1YCf0NJGIX
28BXpI3izRLVKwLtl7zrLsNimnZyzQvF+W/fYFObHtrlgaDX3WZleuefjTHmDVzZ
751syjJL7h3aY9o2Mj90KljB3VjA54RNL9uk5n60XnV+1zQV8TNjl9v+ccVlhW62
7U/jIxqxYDESYWiog53t593ho6X1q42Xtpdigy1c2xRaTE4IJVFG6LjIA/inSxIs
oEAYvZIA+vHE7LUq+hUXH1gmE9Nw5Bx6aqEmA6o6MWbCJ6u0X/Epxl1NMnr0k+pl
4GfsmYpD11pBmjdX4YHSM5Oj0uL3FqXLT6abBao8j/XS/40pu11vKL0zJdR3Jqlo
6F9av15b+qKF8AhWscRotrPdz/sgMhdDcr7PI+CEPbhGDH/1fURXotLQDWN0+eJd
E5m7ls7/bpm0PXRuOCGffYoDL4eQAEWrIBH7z8E1iXrX00gW6OSt78SNoxhOGqjm
lZby7GjkIBKQqTaG95+W9myaQU+gzM8oMd50/EhEeASlRhKB3fXCT23H5cHkO3QP
iFTKVWvYgvLzS9+vRr5hA3d49R0eI6513w810W1zfDehEdfie/8Q2sedUEAhGJGQ
KdH7Qf4Wl3haEkRpNiZ8Jp0QQ/2kEQxbabsKuKhqNDPAbhcEdk3kFAS4LAeM0xfo
1xL8ec7OQ2iH2zSOpKpHzA/eAeYi7aV+B9lhOzhJLlFw2ZXN5tORSETEv55YjZDE
R7ycIz3vyhsocVpnEy6wzulpobRDjmBhs9iRSmxq21z9SPCXBgtUg5na/KgQ5J0X
wiIIH5edyQxJvytK+d/0Xj/OCev6JYTMKNTTzRd0iZe6Fyuh49Ii9qCNQr8H/4mX
Hm0RnIH9+LeqjBXhqKnyczzP/tiyZKdA4/dT9H4XcHMAEE+78oULVuBymc4hcr5R
eVgH2b7OszD+lretautm2P5ofK8U2aizOMnbO3liAF4/0ZyKqwrSQlSXMl1ePLei
DeBOZFXOES7L9w3w3Riqd+dyUtwv0MVpW15KOfXHJZbK/tlWCm3kTZIG1fyzR6DH
fyIwUyt1ctSaV+cixeU+1aYn9LaTn4xfkGPfB+u9jZO78/Cud/gJh7OIfGOlwDBT
0i3aMfQH/myC9WM0Tb3smbQCM/wgrhLSuwxo2O/v2NifBEM3LQuIAAB5ndpNnQZ7
xb0Q4NpyEsjOzWVnm/tpH3gfSHayLIxY/PT/qTrNb2g4Rdg9K8ef++s2Eig43X3V
KnabYOopOsT0bV2tsSpMg05cxEQoDihFkc4uB2QRYGH6Yd/Fy0LKtmFJFZgHa7yk
WCIrp/Wgne5dkM3URAZBKIz24kj+AfgHgTNlpTmHTohnkZ9OKkYe0WxvPllc8QHf
4x2ktuC3GnMlAAIYTixOpBhUeOakyrDGFh1uGgl01ojmq5jHQ1B5P7/ajkADEhFV
1DdxsS0QGwzHQqa5ofusYDaneC0nD4SHiEkUejv9ZooVtxaZ1OmS67ETbGmMe+U5
UEH3Y9Xybqu2MQW0d+07Kd5wbcKve+nxqXIHgxnk+ImjnEBuD/UcOsXZwV0BiET3
NvT14KKu2S4O6kPrhkUyZvPEMm72wQXXOT9+f3/wHaTsj5XiRNOcaOStY+3tqcjG
/9bNP2d+iwhyPDO4/ZgvAiwr2OICISmN8wnPIpNvqSdShY3CqJorJaOVdEakaZIt
Uf0VanjqkM/vjU7OZg7x5RQuX4jCf6L6u/oSYhxPyO/8aDyAvP6nhLlnT+iu+wQK
dd+2DS6av5hq9+QXk1hW0N9rSZvS03nR9amFUuOGSLTRzNR/g0s7hEotQHC9GyIQ
uXP3QZwnN+BSyVGXikng2gyCrs0YlYcLUKthFBhhMm8F9ELyVxpC+WluSSXGFN3c
WI5EQ6YK/P8/PQDRxExJnsHoNt7eLyS30O7GGzQATxTetSj9MBrnS16PfbJ+iSYT
r0ISqydVUR3P83N5osSkJebL4XPw0a97cXJ50jwdKP9ehqJT/VO7EsyYRRPspL1l
ZcQfUJWwtBUTgVRXPhWFHX0jVPdZVA8OY+0qiaceyvYVKHJwI9Pd2qgkXjFu2Ftm
ohdTtMP9A00QdZntwfV4hXrDEE4fFkGBvamlPEXDw3rpGURVFhuO8SbERZgqd2Hk
uLJqklcbLtKSXN3uNfJg1feKoAm2kqHgXzUYeim0pmsdhNbtB/MWaP3lBMPBJ0dz
aMqw3SgYHBswjTBPUXkvLOn93oGxYede5I6f1VsTcFT8ty9id1JUM0QtdfwVQwMU
wK97ndWHkpPdbMDGwz1QSW8JvpLBlNXuCUkQjPwKmBqJHQiI64rzykY41GvCOdhb
AJbQBjUHR6Xp2+wg5tmPZZwBJ70uFp9+OWvcdkfVAw6YdQ3oL3Wvt3Yo163O2p0q
jw3Uk1GeVH22hylaQq5yRPGbmNrdbERWFN98KNki2ixlUAfmCMcKDHFyLtNwal44
c5fDW0lUNQxxHY24RgIyozOFR7OyXaR37+QsFitdFHqo5gTZOFr4VyqocJMnAb2X
2ImIWoFRJgrQpPYUie/I0QWGvSG9UP9SWRWoXf7URsHjk0wXpjdRUZYbRFjjfyvM
8uSglwPcPwDWmGPyaCFMtjrJZBI5JDnDZQ79MdicAosiPs27qayoDJ1HFsWLzj9K
M3Y2InkFjtQ+sVvRZ9wECGqTOtOmAt33A0HyFkysW7ZCnN9x33r+TvRtWwipqB8v
gE/tQXOvKTmFvnHQA58hqkd1YkIJr89JL+DINP1sZpdWiI4ikE/RYoiqHM0cMvGJ
t+Xe+0A5KqYotJVMZ3Dpm+TlWyfte+hDnGlrDygULFrdfKYQM0+omkK4gaavatLR
U4aoBalDhb6CEnssZ6TcKxuaSOgWlAFiTEDVCtPypOiu96MpvvJOT35ZR/i/Nr9d
FkngOZ+sxj0iDInaVsJizJnu7/0oWWi+KBZOt452A3gOlJpHMAr4oB5Ead0wWvU8
a+QB+AxTgWqfepYs7UJETexziEhf2ZJocK/99Ccdx4u1zUzlx0S9GzC3t0wmewbk
7CoB5dWEmHKHyz91T/NYJzasxiUzockd+h62Zu9zvfe16nj44AwN3IAdu9EZKGUA
TF4iJNsFQRCboGfUhz/gL5GDOZldVTm2MwLoSFBer8HhqnK8pefEXnqFPCuYBYqa
VTUUQlV6OIS+VB0QnvxeDn+i60pDq1gIsznTgr/6kHMh8OCqWr4eOKjbDqKQTXgE
MR2t+lQkXjATjE5yVnZ0ESngZERSRG7RCNk6fMv06sPmG/NfTS890xUc5JYk3Vme
cptYePCzSeAERgSmUok9iXlqDhDC36U3yn+VsxXy2HJugGFWwXXDB3VOnVjTYSsF
zRFFTrul36bEVeQtSOwwz2gwtBOKz1aLmw0S5uJQDzLRIl39fVaj7CWQT6HvINRJ
N0Eb8Y/yi0lqCH9y/Q8pNgz63eHh5xRliE16a/dNYyvw/j4v1B0SiBonbmOSXlgD
B0szDTYENsr7/ZGAwwCaB0ppAM/X4TH52YwZxzPeW3mi31s6c+WjEhkJYyyrW+tk
vJKz6WlqBT+d+A8Af7TOmmijEYoQZeqv6FxEmTQrjzL1AcQo9Kj072/LV6h4CyHw
0e2ZoL70LvbsfFYLAYjW8a/DzvGcARR4gSsDFprL9qM+GDjuTY9FSovfqBkLYCA8
y6NHwLge3UhrIhQrI2M6LbiAq+AnLdbS73cMOW8YVlhNiF2iaM3g3VaPxnVNEGat
uFvI28IhboC9NbCRedlSRT4W+OYwgsKsNCBQQbskgmvNMbyo5IDGOj0FL8XEzTol
9WN9Q+9Tiaq5jFijWq4Js9SIoFzFanKtz3bT3IoK0HKdcCgN7JSuX3vh1s3C4o3O
r9/bdqGWY2xsGTapGdCNfqGJeMVwyjf/noeyJETZ2QjuLLWCKzpaUKhU0uC7PnYZ
LQBhqQKi+eSqQfFBnhb/KmWIsAS3mSjfI/aWo+/aaKiHwlxbNiP5BK0DqqB7U2gu
bbzymqVmS1FmJls/GeieDyRtZAnRQPAtpfMDBl2Owb5ONZXuAjGKdMv/5P/FtwBY
HJW1IpFbqdtHhcD1s7jOuQgX1e6y77O5Sc/FS8TeKT+M8CJY/s641AHoMpi94E+p
xxd7VbkzCKrBZRfqCuOMCyAxqiNxd8MdVT4K/Ov5/ENe4VsAN47OSf4kwMNWm+MO
A8zQYMChzxA2NZE50ds8pR6paXyYF9/I8SCidmjNQGC93o3xIPq45BzYJWZk/w1i
dGA1DOpmJpV2re7bReHN85FRQT2Gv3DCsCb2RuE+33HJuJLohubedkum4DtoSkyx
5UkRELelUWzzKt9h2Fi71z+WSPm5bRh0B9JSjGkbktDQJP0pZdTrl7ZRAVrZ75ST
gTTpTO/5URH9loQCEgGRy+ikv+9b/TrcNCn0wDqk1Tq0/fS/yYQYd3FUJX+P207Q
+/vWlp2m2p/t6H2IgPwVezBjfkDFiZGHPTtTSStCAWun9M4B74FCajrdswWx6s7E
Sfa1RjTiT7b/UhV/Mhg6w7xqbldFW9/7rC/e0/VNIOF7ENnbxtfyHjHa/uPf1GKn
S3cQFhe5CeKSYLzzKnGixttSdUA1NX8IUZgtrdmii+VwolmYaYlL0UYJ0t1YpvSN
JX2e4P7ky6XVZKrtTuBeY7oSrB25bib/rPfHI5HiiZR9e3xl/b0cbeq8/CoZ1plX
is79s7lNoCHKsF6DBDKD7bDbuxs/DUrrSwubciu7ff874scOsTyGxYtzoajWTJJp
UT5UgA5eOxQO+Siet0YgdKdufBynq+EmF4H4vly8ZUxpPj9j447XeruVt+b7kZ8q
NgU2TvEEJladNR/VA2QMAxhjLiW730neszJU5DgW/lCA/rqD9cJg+Baku1P2zEjS
SpmX++8eAu6tZLBJEWiw9+bHqgLP8HtHd8Lm/cXQP6Ejte0KJuSk8KRYpAKhFd4R
Gyg99xwPm0IDnLYCCemaE09g/8vimONhbMW2E5GMRuracTJ5CG1ccyC2r7nSE8b+
4ko0b3aVeB0pi0hYr9IKEpzN1H70v+u8HOhQu/gBhnaANTZ/PhuBo/yjHZwVW+m1
EXjqIi8viov/pQx1JjqvxJGnoUuiHfbA4vu3pPy4quT70R+7JwGZSMr9pmEqNfv7
qO4TjBdDQiCCRPkOmkQuUWbiUiY+M+P60e43QOk1yN5X7ZVdhN3BA2s+qF6z1jVQ
lDPTcAWJjJCCocNJnuPd7fF0fBqLJpdYGZHIg+j91QxtjfUTC1WtG51hrVPt4y5P
QHzOTXp+4uU7V07fbayHBe59X8JHRByM3ogavBBEhT5sxUDiWDNYIiS63N5L+98m
F9apOGbhr6h21tGaVUIRItiMV+qu0I9KPb6bOi6/Kte5jfD9dd12lRYW4D5vu8GP
ihU5rcGp/yl6EDHDlI+50hKRTwaocJxuAxry8Dyc4f68Jp9Z5N34lSaMdrp+cfTg
OK//At8P7hOg09DM/0jnBnLfktmRVKwDW77N73Tvs+5IImueSWA47casWEKma7bC
f9blUZ026DZDataDlNJjPbAB12thVJ4K+A1eh2ZdfHVbzjZ+eowSNhFvrPvZ5uiX
11jXFZwOYcOzn7YzpYzugkXdbD495wlCNKxJXC+JwuoEjOe2LwyJHCcHyF3z+7nO
QhOnv26AreS9F7oVBpvGFa3tbY/+DjI4OxV1r9boDgU2j4FJihyKa724x1l1uDQd
pioup5CLCwRLzdlMH8knoiSepn1R3PwZtVd9bT0rcH8ao74Lgx5vf0f+3DmQIMda
uXpV/z0q9eRsK6P4yj5fPTh2EIsHkXQeRrCpsGQcMeIo8M91WLvz85EndrXV56FM
TNqX+UeEBGTNoUBwAthGpn3vuTX06nAGjoG6LrPhqa3PD95GnNCSrVaUt4ADdpmV
SNCS/8DjQXeGPIk2AMheYVrIEV7iVB07KWnz3n1iXjJ/bPw/XuPxd/sqbVwWEllj
DWHG8aphawjkIfh6AP8wVhIy5+wY7M5hb+/wmZK7T9whvgzZhpbO7kI5zJHcFGNI
ySHXjIVAdSKDsUD10wQmWkKEg3PyaCKxLdpb7zoe5bVSJBG9czmdkLCu3lAwugeq
iNfubQYpp3MrSmOrPcZeOS304Jsd0bi+Cqj/zOnM7Zv4dPgSh0PEc71MYkZp473l
aR0JCSNy/eUFe7yuln19itqczpqDu/thKloPMQzZDns+ViH7XeOAKOwGjccUO955
yMqu+1F7n2/t2J+SZfitff6MN63V5/03VS9x80lCJAfSrwVAvxM2B5sHGwseR1Vm
5XIoDDJWBTWnvzu1lFqQENMm283tKXv0ioCfjCLVjs7MnbepNQ9X32fy5p0jF6a9
jY6HM5oFGTUAQUPBF66LCCo9vGC+jQf5pcLOFHtfCBPfw/0Ed6HPrBJ4BoxPcMiP
5duK7FA/uuCgcGYc2tQW4N4g5FOdoRAwsu2AETR+uQA5Ej45US7kZn34On4FZsb8
SAiqQmvgYpftWxDCC1XsEFvR4GNawJJGX51sPQu3GgW/9spk+lOD7WPUsCceURrI
8YrA+mj0UL8la3eVjnSVE6R9HBI/8wMM1CZ3z9RW8A9Tn+5BaNBz03otSKSKpgI5
aBwAzoRZVE2GvJGQNGcwpLmFemi+fGEaELHLx5EJEOQqwai24TB+1vcDb8gNVzEX
badoW96Wu9Ie3h5QOPTpAI2Qv60vHXutvfdg01Z76KaGHzX2w6h9FZlJCBU9b/S0
wurlUtPrubSvEyvIRzgSoAO1WbEuWJizSthN7hNNTNp1UX4vb0nF020o1/ef0S0Q
WjVO4PIhPBjWz29IlLetuoN9oDTEm+7C2gMFu9D8q8rt6rLuS8te2FXPcgCQltTX
cBpgL31U9VdR7/ywsTLqxy3wRB93NXpNewMf3uQA8RlsDuBi1+5M7ofix9nrLd7a
bZimyuGi09gW08GpkdoGW8L2c7kFupNyvT0Bu6KXuoAQIMx4Ax0f7WFMse2QjUs9
/BbOAx7V/A6f0NMDPJzmC106pD2kVRuAN9gUAtk/56e+BhUEnAO8pE+fFK1yD5gQ
UJvDGWVLm9J77h4+viVEU88ENle40ER0zV5fS1FHdjQDxQvC7nAtSpHDciI0J9FV
G9rx1DzwHrILAzZuzcZGlwcmfhfDTNStwXoW44n2P++N+eANKKuv993uc3Ou1qmt
VsSfsfxT1KS1v6qnl8kB7rjpLx301kHlhI9tUzzCJRD5E1TPUAFc+AnfEXJ6H9sN
A3S9wh7Re4OPI9Qbub+ahsppPU9BPVEMqm+q1AIG+OXEKA6slWNKm50/5FbWC+cV
+MeWcQOh3lL3mQ/dUhyccyvLxkQljZO85QVDXwBuaUAhbAdLBysdDCwmuHaJ81B6
AN0ZHKL6ehJbS2W1HPCSkdAkl7FmR4hEFsZSpe76hv6h50IkprtNkIfOxY5IJG4N
zSIxCh/lMajYS8i+fKEpzjF9Pl1tB7Tb0rMqeOVCyT9PTMjIGT7z0Gkc7yt/ZR+3
0vidVB0AOjsojZjtGDE2bMJLb5failaoTNzXa4hSwF7NgwMl3vJ0iLhqFihsksDA
tECwYYNvYxzd1cLZmhJW9conNVXhXgN6gPgEHH0ao0+BOur8P3qRQGsVSj0Vgiqu
GjW45Xd+PSqSVuylAuziNgwOhJEb0/BhbZmqV+m4jv9Rv1M2oa4O4cYK9vibZHRc
N7trBBZU+pFCnYPa3hCgie8jJvv2nKNfKgR7DZYeafFpX6N5bJA4Bji1ziRvEEU4
lmBwVwdSray+XwLyGM86+LezUeeKbtyg7RtK5v8BzhFAsloU+NOmXYXftniwsCYD
yraSua8GMi6TNk/N+ChfVEfgsZYFba8m8uNnE9OReXlRIV4KEmOF0swGXrgU5rON
hesTgjzUAv9dyPO+Gl8zn6Pg99CjaMwLRLWcDsCTuDD6F8klGFwUqIsEVKI8kMO8
XYiBM3GP62vu3Os9PHRz7UnOW8jMvb9RgCO3iM5RC97OG7ukjFxb/FA+WJdIPgin
70vKnAvm7h2Ry2YLYphSjgIit30ThiI+juyTGklEaL/R5s1W/bmyi7+dHPMvcqiB
cj4W43+enmp4zhTJf3qayGvYZQ6JRadekuyIoXtOpP0t3Fde70RZ7ems9IrmPspp
gU46Eb0x4KiGBq8asW1dVg==
`pragma protect end_protected
