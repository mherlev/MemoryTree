// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:52 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
RAIdqL3gXoUO3ytFNA9iLaltjIK6/Lg/YQEopXNFCHCQdepkLYqbk/QB6idvbpub
N0SH/hoXWfOWtcR/pxnK0XOxmextNvUd0pWSr3MK3JQGbcmXqh/CuQQBI4q5PvMi
wCwhJ/u/e9REN9uxcoweaypHcWM10rU4hY2KX/N4o3I=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19360)
VBiGIIhe4rZzVuLsCiEM/+EAE/VrEZwQz7OpquWAxDPTbFSeo8pJIlXHdGK3jOip
FMyG8vaT95YGol4nQW7tBvTFLSFHgIXWWXVycOjoJiIdVwV1kwvu+njLjOtbhY2k
G+JVCN3Pqk8xr2c12P1fPVg5HxwyGMeqWf7kTddbVSqiSYF50EIjtzGUf5+DEfqG
24ctnnlT5Kq5JdMAFZZcWkhhAbI9FILbG4IOzoxxqOOx7msNe5BZ0tjANZ+chiiK
z0oFnlSqbCP/Ox/wnPFwdoQF+5wqYuE/UQT+H2pB1on8Yeu0bvI2lZaj/GBVdNnc
a44x/HsQjQtGAzdgs3lm0T525VLqtM1b+HVzd0SwgdHyaQ8kkY4EFkkoJvUSt/Uh
1nQnAxcwJLcZvK30EK97GMMc3vZ8o/3TuVfblxhcf0wc0OaDvdMmUcC9PKXNDMuQ
xMctyxzohdUJvYPpvDJ2nSdSy67O+bY3pdqWXzlhTYqW+/yAmcaoHDrDqSXIzQMp
z7TDcJ1cn+m+tHIYXft/T5bW01za8tV5Ud+oBDyCS8pPkdWe4hYOsWKqRcpXDI9z
guI7nSAeMQ63BDFw0zBNEqreVBfqVErFqs1ZN6jrQaOFljsHCOP8YC3Ln+m+DUD+
0/SsmEi86X7G0hnG/GufCjkfy+jHkPgvfLbs5pvl7vN/ZOGjrBY0g9QOwsx47t/I
g7SpyyyJJ1rtJ1h/0DlBcsSoL6o21+SiaC6LdurLuCwC5uMDykHDpEFabxTtx05d
fWwVgFznn394a/6t+6ilOfg1i7AIhTvsN/m4+iuojxtLCqJfDhqQrmREtZfwQTok
/YS8hqVTm4h72EcAhoF3nyJv8iEwhDx+ND9N8TB44nk0itkNci0AeI+nfmypY7pt
tSgXZ8KIVLvJM9kqCglwu1c9qxCpdHYjgxobJQ/wifpkwveTpbmDSSJXX3BfWHNl
3bfpVX8OVIUlealT7netx3vt8H1cJzCm5UXx5Wb1y5qEynbOKIKAUDjngoRkgdJn
OTlHrhfZUQPEqpeOZtQ9aTCMR8xoBnaYzfWW5t6oP6w9jFO7EpYFeOERH40Z1l9Y
E+nKIEAHY96smw0dOg1MjlhMBM4TEiAFSSAvZPJK+m1aOQFFbjiQM7deJFHGBshZ
48YFwksQ5C0g6nGEQiNsmuwt5rzov7dR7Kz0aHOZjFYEbqoPlns2u5I8xbaqulm4
sIXJpMQ/MWFzancGRU5pV3Ma7TXX9f3WyJnPOYYDAc3ln8C/j+mjQrFLBOuAoTj8
7GrH0LqbfB8FZDO+pZ4K8T638yuSAMfqdntZxfSS5GCs7c7L+KHH0iO9N5QBLuiJ
u4cL0zSmISqoanqEoYHyZrwK9g+gsJaB52ZAYPG9g7/yxXW2RgwS0KYGAd3XGGaS
KK9PxYjY4D1lgIJtBG+V4G14yF6DftTD17aK8ztiKJ0sbyQ19qyzNRZR4eMpmnMd
bCvzhed4+45OzKJhrvUIkwnH10GbyMr5yA4LyKvbk2uvaWcaqdghWQlOcdJaELRK
KcGXbRGpVx3gwyRw4C9pPnKX4cE8334lQeBwY/5t+ik+d0iaaUQHQdo8cSaGKmdN
FXwEOffv+gfGTDe9f2vSLkz/WImKh455zMzogF+kIY6/6cWDSy4hfNfIULoPhoTj
DfiuNaYXJ6iR1K6iM8Qgor6daSOVw43I/wNDbBcPueQb4dkqTdIs018PQXZKP9Qh
ryNF0aNpnZ0FBMQgiz9Xd7QKnb23Rcqul8hBi4QsyMIKdEOdKz/9TAHJw55b7ah1
e9+ujAgZ8iboEuUfIfMIdqwULinf0qp3F7tyFRgZPXv+O6CEDemRVln882LwkXfl
/ABB8GJxi4smDl8yQ/anadcbbSvAli7gVhNg3rJz/v8ofz5mj/XmgzDcg3tOim0z
ziny1acEiKTwQmCKO8R1HzLgIH/XMNamotKAuCWXt2R3eevdkI73oNOS187mY0w2
lG4a4g8oIeOFuQMrsHZjbdmrWTOenky3AoOQNhMKyHAKMgGcquh3m+SLDEqxLY6F
JRyL5ZPusRIV2T+VdcS38eU53Uld/L6ou4XXtcFB84xIN/JTV3BpNr4JwqdczwFI
/O3zjCdPkOxLYqPKrzzHx7NYw0Z2OFxa5vaV6q7suR5edcSeNbandoVUKTnS803i
mKqihxOEwNqufh36a+08js/BVqMd8Dj6/sZbiuYBB4xOTdGwDWrZ+tbJs4Lod1Ev
bMT91HazJCmc/8l5Znt4h6quX7nwsM1nycxCx/enfPExCj3QzoMODEzFEoNC+Fae
EEgLBfdhAXQjUm5lL7O1oCjwTYcclppUOEuUuCL4S3c8KZDL1ejxBWrI3eQHbNH2
WdWM7KDR/nBdg65UhS3s7Aod33x531gWEwj47OHUj0Qh50rDMP6wNZqzOmj95KTx
IcL/b6CaTMJzfsfK5gmSa7xbpqKB/jq3bI1/eavr1cRdZmO5F0CTSbbLZ7+eAvgu
2+TFHRsmv6RRKRhjnp6QlYswcr2iMTyvZxAja179LoWFlnpjMOjCxL2VvOakkTIE
M9vcaGlFLChNgxbafunTn5bPH2nDb52WWUVOXbD6vtNeqvfVIT1JWcaCfwoKhkBU
+y5bXwvYYlspK/QfbEoNggHWeSws6McSHA+eB4KZCIuS8LFwg5sNZrfpdpJPIgqE
orOM5130L0uFxKLYVbWqxRP3xe5+O7R5uU4MNINIVe5ZqrNMveLpSeMyiP0VPxaD
SPiMd4xhr5LKx86W+hYSe2x+G7IO49phCgOaHBtmIGn2jqzSQEdEvwtV1ioW1qzU
j9ZR0MOHPtei/2DC3tJJK2g7xd7PylXYlx1VDIjuRKdxfWanSgYQem6Xo73ZCDBg
JZ/AXsJg5bd8EdISk/NH0PcJw5c3KGQudoBhQJBGH3Nbrk9U6yrTiZLUCgxQPerQ
Sc3+XkKRX5+9nb6j/wjaJlmVCuLUasoER6PCLAeJkz4toAdcbAePS0vrJtPaYY0F
ua6thJb2LYTzvYfaxiaM4/BOTfLhQdmVQRE4vS7atGh0M8Wvs6HmxXtugFoTxjkL
oJYYZUCGcrUJ8vZxk1qT3EMVn1CuP/x3MHWB0zE9EqRnBms52L3gvmGqPGmecupn
pioJ+GR2atEY3JwtMCXCBPBF4y+xcstwhdgrlBSQ+PrncKXpGfFaIesoqG8WEhrc
aXGNGATfkrZEM1CTtsjNVlRgrh65l3L9qXTgwCgwGJp96r+G8hKX4/T2ca+SiltS
cqc7S5vTTz0M2JCB5BKdh2Hrb1xmP+//sNPDLaGthg0JsDHjO6a88kC6CgRgPUlC
yqZ3WHMwfW15wl+rfgcHj8xlqVx2mpDN8c5JLoCVS2eQyaddPAgFB5l0sY3Pn6TY
VF9cxE5lPNYsswm9MYhc3/7MMTv2A/BSI+e3zD6ASoNKhWynFwDu8czE6WTFR/+O
IlG/dbpxcxMqP8OTgR+l+M5N0nPDwHjX679Mx3/pUSK/ojJe/OAGCkKxE9Sik/5w
Rpw2KRi2KxEKg/XbQsPfd2XYKuy+ljH6+V+3qX+0WYJgKXnvlDgcw58S8hVAtA4r
1InhdxMvHCdnvlOzwLByTr/g2nKKBiJ7xeR3N7YK8byIes94hcReKvW96mM8/tSS
Ex3UUMYZfpzcMhuGPXfmo7w2FY0mLhe6hcF50YBw+4LK+PHweb08B/hnA0SpOP4r
YjpaKg/Mhz1o0fKz4Ic/Vyk/H330ZwP50wRBKfWFPnMmXQQMsmP/bHpjXD4l/qTA
KLhs9wNTCiGvD3LYo6y1f3sOxqhbhYOyWIWI7RxDT/F+CprdARnSdHqlT+/kJz0L
CpvU7o+1tx925q3E6T+mylIIyeKSDlUk1K58T2VtqXSoSf3dG765XSOjR9qcEXOy
fzoTZkqoTR6rKXd3uaI9KyrUnLcqCJPyNbgp44NXCFoSznpasIP9T9T72pd1DEZL
YeU4aoC3/V4/JxnwIgEIWhgdeaS9xVaaKOkeT4/1/T2SEU2VTkia4QHCXd+V+W+8
XNeZuyovdT//h7uj+XmGv38c+4C7YGsvr1RKIWXUtuylgs2VrVzBrQMhdWJHNHeS
wEIDuOckwBZxvOctrqXU5AKM1T5vS42aU8lItkGt8/HR6SGaeC7jZqMvHuoIDiZr
qgniFxMtBkihCVNOLd0puN3sZVXkp9k9U/GphLKSYKMmZm9tKEFPC4k91bMlYnWZ
J7ACNh+LzGyo2V103NzzldyD0j2fdyOJnM10Aiep2b1HPUeOqi/itLk10Wgz8AzU
ApHeqVX9h/hzQUIzVqRnLHCL66uyodXHDpCubMgOmmfwDku5N2UhE/60QBNmwX6s
n+nKHMvq6zjUuQlm0qI7lnHiRMiHfIGm+sYXWhrGIen494vtTdLZHEWH1yjRQypU
Y492IVRTYEYCoc4Acc7Ht0kRsHlPzGjtm6cyk7h8RccsSDaqxXeiTIFo0+LszF/S
ij6DgKCPe25E6hGwxw71r5LaOMwtWw4LlzP2DnbLI96ziT1cf+Hk5eAMntp/fSgp
2vPLlcfw/4i4xaePENInQnQmhZfkpjUvwuWdayNMLUvLvqJMSQ6X/FDs/4R2m/Zg
Nn7BnvzCN1bXbEQqwDGCTWyRDr9SY/kY2dSaSPVYx1ZUo2E1U+qSMvkbs0ziktjn
VSm9YUiEYoFZYAFR6Hjb5ihfgVWZdXdErAanNzuIuJDSABP83I7FYayRS5e5x4jG
NXfZCtmrTxbTumD0sReBnGKPKNMYPFfJh4vSVi+wQHdf+sawJxSPYcp/Lmi/szF9
WZg1o5dexZwtvVk3gmMTljgsmY1rvb1vXiyxGMINFxPZkb9+xP/UlCkjJipMLL/e
xI982XH4o92tehrARcFyip/cCZALRliXpYp3Q65iFrU2ttP0/QoCyqmTp25LWrmG
imp8ju70NyVD6LJuHWOcAMRDeCvo42mHCW0RpvqE13JdPStLDTRsVrjGD/7BXbFv
43n6T4Uxn4mShgtjYWpXGLumd7ZuhxEruA2d7lSsU7daTcqhy2f0OVp3B5fjBhY3
0p9UHn6mXsccDeYpV/2pBvgOO7el97/NmcFwvyejnL0iGL+1/cTatKktWA6fmKVX
LHny5brB9EfF9RhJJFuC5N4BGs+ZjilPXgdPVCUZvGff5WqISffTCCnknKbhdivP
QBKEPAu0Xe0KjbFuZb3lnwcItYfk1JyGIqUjCRrRS/82VnNjl3LCoEaK9luC6n/1
IZMFyivch4DRpxDip4VZdRBZuPhMk1DfLq1DktRXeKq8XwjZTsDCkAHHMy43jhpG
oMBEnSrHYl6djKmLaPn42grML16tg5jvYB6MELCev5Cyoe7cdZd10z5nfdZW1ZCE
9ySAAbxInw7TS5ScwuzylTWIhz03siKq9H4QtB7pm3XTOwlupsmLQZ8U8fUMWHMT
79/4/CXrf0S7gOGi8c8Q7/P7W7+YbtKA8WwTZMeLC/mEXP6UKxmcjFlZm+DV0nrG
EZgtNz45ZTILmuSQnvCWWGW7ETIV925JDgwTqIyGJMeG2/t+ondjwr1jh5WJryhT
1AymM0oqqJ11F+xirxg4VRPfxoqCc28AYwNKgE50XnDecqMy46LnA5KoRyrx6COB
Yh7uy6+hEvwTkdhdDznrHl4wyRGr7M06zzfz9n/CLhWGKff1wT/evUt3bbiFjb2r
bktpGMvTf6GB3laMfbcw5mGsiFq99txZ/f6vyN1eUmvgsyO9ZSe+2zuEVk0sQMIn
BIf+L9IVq6Pv97vuon2CFsCVB9Q427eUak9g7rtoD6Z5VJPMiLNTD9IczzShUeDH
yNlaz/3rafsErHwhfVqU8Y20d12Gmv/IJXtUNPCQLph64azarTBFgzidbqQa+h4/
gQdBi1qotK+uksba0L+d5+Y4eyZFTEJerMwGA5AIuasoFWvMNpHi6S6wSm9uzjl/
ryU/sWjnRT3SEeKwoBIW0a7nqYoHLewylMTrCcRL5BHQip7bp5nd2ibQM11FUXw0
rCs0MNtUdruG9ywWYkCUS5XOWM2ZvxwN9HDaeYgDtWipRwkhDKL8Jr4/iz0Bw05P
DBEAEDgGBRqrFWfZ2GcVHW51e6yYpOVb2zGAWKgbC6xbJ/jYIOGs4sJt+ACyu0gg
T+ZW9l4nNKSjP4D9DjgqJvpmjyMn+0g0HItYzTt+PnwQETVzH3g72VYUGdWKWxxw
rcAAEIoKSGJtXUWRknb36H11/k3zI1cCUp70S4vjBGo5VgGIXNrfRYK/74S53qKH
JAFya+HzwErLzeqow70XT31CunKC3unLssxbN1pVZaVIy77fwBzWAE2DBY76F603
s0Z0zj++e8+IR6wfSb3Iy/s6bUSHGSv12fYC0Y255oCvZkeIWWfb+Pqusi928kmB
FhBcNFCV5BjDErbGAzzAxCkvLkgEJ/yQLj+G4i4m90frjOt8orbLYbWqdAQcutab
y8y5tOgWw+8f2RrWSe6OJIsuo+26fR+WfVCnb3COrifwoR8Sw7JIXzLmD+CkHS7i
WROVV29LrZupIIi1qdMyHiJVZwECCAtDg1SOTXroCKO1Yvc64c3dsXiQvZQVprZ6
lSY/smDPDcykdWHIvBm9RALysH9q9Hr60J3mGwwVu7gILcF8ofTn6M0rY0L7E8He
AexTu5LAP+/Ze8s3fNxVpSA/+rTTSegYFtG+H0Kujg0xvbDhlDSGOC5Op8seCm3o
W58zw+5TTjUhCB9hMNxgTlelBEnbpDf9I/zuGpmVhktqo9dw429AoEt8y9vmYc8h
DZwpvCS04bUUwKgLuViInMegOJN5kII14lJf2zdDhzKFwQg3VA5b3lfeoe3Gk6M4
nUZ7+A9ApZMVg+EmEwD5WYjIgM1X0C4Y9c/t+IczNWaL/oARsBjco7vtEzadKey5
1smsd0HkERTyRLY67rl+lUJnmkUrJXBDHqfTAACr6dXsIxDdo5465+CoJ/JpIO7b
9/H7ISjqNv2K+bJRRj1YOE9Yg65WU1czs6WLBqr4QnziaE3lxNtr3VLVG05cAKt9
8QGr/TanrehugV4K+TGfndD/XY7uPusV7wzOBhG3igXNMLz/2IPt/v7f3YNu5n8P
Rf/Z9V0ScQUyFF6evlnRtULaWcJCgo3xCt9G+Z0ep4SAkT3/gq4b7UafhX6qDN48
0D5Qjq2nM4lWcIRn5adoJtXYXqaDKaCTRxzvYE6Ndy0zdOsuZQ33jslAUiN0AYyR
uERIQEbgacsnG2BmUGoAgljWq/lyaT12pK7mjegAzNwRx8cpaHTmfpAtsBTBZfv7
vlBk+JIQnsRqUBa2NZ8khLGQPK89TW7Rbo/GRifFyDrVVEHIsT2EbX5AINXybEgX
q9iLMjUYIfX1HawzcuicVdAZoL3sjX10KmeirzAdpoSXuw3OF7m9zWa4xFetyW1d
670ZXVwZXgwYjsS/v0l+losgrbLl1FEO/I9+tqgHdnNT7RJABscDng+hr1UoZn2B
E/U9grCbw0yOmnhH/5/QDjzc4Keiwo0lgsLIplGHuRl6znChy8+DiKDx5G5uitJ1
staBBfE0CgUaxMDfddN3noUJIQhsGONk4hJb1D1sL0Jf5M8Rykndr8T4W9+Y84Rq
cav99ywBj6EWxosaUK78JQovCs5I+pju29x12dcUgT11GjuEW+rT6kBbckhPERvv
hj2WrMt9g2LCtuwgPA4D7dl/0htzzwbgVHAo51VSswAI9qdSOe8hnuuSQ90UH2gY
AdOLQ3aupNANmypPIjzxBt1ks940HQzv0kCJk4GhT3f1Ys2pArKRQnKG3VlsFICs
3pu1eKU4xrOVC23ZIBc1dix7UHJ95XB4gr/TzOO5kRNG4Cp4nn6yXzQClSMsRhH4
OWDDgmCyu9NwxIaQiaiTYfpe65UCR5bQpieu+S9u6FlGvh+3j1nnCILUCtjr5rsp
MciUWKK/eEU/4AdV1SrZRDmiKWgqWNJXGodjZMweL7NtnF90xpfho7sRvSj/r1V7
VhQn9mocsMtxc8HKPdfGaA91iExdrxuvCvwLfqRb73fTyyggqmtQbKmCwXSr63TC
9HDyqWL1EPo0z/ubQX8PMlbQLyBeYG3iZ4Qry3qVDLZLmW9Kk+EgR5hw9d7vyUAg
Ury2FTJKld2Cbpl86fAoheM9/ZeJpPkehwIerIzyQxs8qQCGyom8sto1Pypz1Iru
LJ03ZC/3JWkeYaCtdv3FMWV5i1lY0AgHm6vhvvnQc4Ke9m0bVPqmVkyQpfXPxVLd
ms8el6vaH3/VmdgGkPSTJqPNNEBnTvUmH9a6bzpAarR2newAAYLSHvQEC5O5TphM
kfG0DgC9i1iFMnZk7U3NEDIxjnFMmqqBwJgYEVPR6DQ5dDO5unix9zNy/xrydGmG
4VZFeps++JA15BtfxxiGUkD0jDG2ASWuBHmH3JAL/34ViLXgiI5CmJLum3gWXjqs
ocse4+SaQ2Up9wne/7VZAeM8799xsnjO7QifPGHLBDVVkpDUPBJWoM2F6mhv3nqf
VfzfG0cxTbD6sl64J7S9XFrWW6OzGNlyYPqG8Wv9fXREo1batMVAxBox6b6S8Xl3
G3GL4SI/Yb3pLEioGJKy/Lu+R93U9q6JqAWQGHrJI1QqgPkzqjr75orosgjgqIHC
HT0SypjEc8lhCoWkmpJYd3ObC+Ff/M4RWduGLNei2uzhlycNrhZAKvKdfnu9Yjuv
AGxWKWeM/I5VWAUtw7MT+ZqgjKFtA11Kg3IxQ/kWoDDIZfb6dujyASMjtD18LrS0
sTMJul1mavNM2n4bL3dAIvYJ9f9+8NmCP2nFTWCYD8+y2VTmbg1GsWhcaAs36L+Q
cDqod6BBNIoUXdWQNDO6MbVn4Z2SnC4U+nlOXnYn+yEdA2q3UrF8ENG952A0kEIc
jb9QCdYNzLA46J2uoKkZPtBMVVhhVS8cApkB0LOrFC6SaplhonL78/myY0DrE3cl
aBKALhRLWxzJZzZpvCU68EN5ZvovdhAntY3h/PAPpzr9A/DqWNkvp1OGvKeZlODA
ni1Vsl0zqCDoG0BxmmyMEtDPMHQJZ4dEs++1SxRNCOvnSEfZ3K22mAvKJhUXX5Oz
gy9wKsG7qInG2mo7+894QJyCnh0/lMPruCVOqtAdy+MVRbWbQ26yooatGJ6lEeDG
xTAjyJRQQFLmP2FRmuC50FpMUyu12Kphx93Kq4gWZzVj6XdJcwFUUFNFqysyJWFj
4qFQf5PIFCWvOKkTdb0HliXzewiHqDyMIFUyBo7KR301q4LHYYHo6l9XxtGldubR
LZd81cOwsgkumelrrjTmMUM1K2Pcu8eduBtRP2AvvPolgHiSSt/dNdvpWiVq4Tjd
zWhse8M/Sk33kOmk59c8xEVPKzNmHQLYEKqsnVWU1uI42nGpTtBQ4ND50De1wScJ
K/1eQoNfq/sqrCaX+RG0tt3tFlGhEDMO130hJVUkHZpyYbUIkqJPmA3Vz4lZdIOI
iHttGP7EqwmOhUE1ObWPhXhFAM8HYbUgrWH5+gn+Ginc79pI0cVtig4mKDJ5rcxG
5xf4avxcZKIbgecUICra5KSmfsOMSN0cZFT4Q+kjmpSm19OYDvtWkc2oZ2uKZl3W
9a7yJ7g8YwljZx1+MJeenuloPCUZ6wokq17UXLyZa23nBHk92FQxFBF6pjT9Le8t
x5OUN40Zat22LuuqjVcSC4xKR/cCCo0EWVBR/zQXEt0SzTxc6s56Mw7NhRPTY3nK
A9Gh5cGjHKVBGuXvm+ednorFdjglinViOgNei+eesY39TWAKzVCLx5dhI5Rg4164
/UrbWEwtAbswoou1Flhu93MpeGmTQb2+E2umBTf9eOsPd8uG5ED6/nqfGxP0nwMX
UJ5NTkK4fypQ8jwjg9va+/LYpAW8681lKQ+qTT5sEz19kpc2BAdA8CxcX974b7gR
V36nUKtmvcJw8YyKIn7ZzzFdFQgvwEY0MH+LKuzxtD7xdEKqqZBA9YA8DL/uaDuz
+ZrdfMOlFBtzTRfnEGWY3Sj6nIYy/ylQF1RTWrmHlXk4kHKh7Z8iMzjvrhcvjkOz
LXKw/NsrK6WSrF7IwNPCxGysnR+BFP53J+xvY0oxn9532CD1xHWQRPsmo8pBREWt
XmTxA0HH6UXXjHrWT2DyeMeGTTwiitTLq+uM/JQ4HYq/udAiK/oxIRVoKTrptQoT
vL+hp11k1WCaH389MstJXHarvg50U0HCuG5kD+cX0HKoHMNgSfWL9VLgglbl+URk
qb8+GYN9DaV352FdClWZiuyvlpJhZH+sc721JfUI/eyaKYjzQa1QbC9u4E6yX2CF
CNTs/W0rftfVOF1QgOJ8QXoCAl5+To+GmpKcBGnP0r5c5ZVmGKEcfqucaHfLKftR
9dPa5v5KW4JzqEUSaT6hoosBFUFhfxe9ChFVBDVUjdiso4rmS3mG7v8akgJsPo2f
8mdY9zEQBOHnGWjAj54TQ0qW0JpK8XHxSDPJga5ECgZTf1njtRRB0w5WwfVqBmvd
Un8MShc8kBkCZx3eRVg8V/Q9CxH75DL2FWRfYJoYkmkGFMWy311vLWfTKKbwSr0s
wROC9PEdgIz0DRpLOXwB6TU10xigYigPEemCppY0Xx4/Y1OdRFvBizswAnOaB3ZK
qTN/UUwM4mxQgN5bLGG7H+nlo4/8SvxtH0ihzzbttaMVrMPKxQ8GvaKhAZOoj2ia
wyozDPDKLyKp/DdPwb1HDEhtXPnP5ZyQiR+PI46n+RMQHBv/0VoVRccNi/n/1FCq
MB/gY5NUaj0/dWe6JXHT+Y8c5L72qZxKXsMiaYeGOYffMvSRKTuAJwrPTFAzHDMM
NCPWUlG7oi/ot0ONBoyQzHUYwLLztCno20BiqZLvi5MSVGlqq/WJb8KNZTJeJQeN
PtvDXPtIbTVYjrn3+96Sd3SAU/UhU5jSNxqJCrk/ruJv4z3sjeKv7XRcT2uVzYsE
xGn2OXBED9wb+j+xQCmODFDn1eyA5gnGCor6vZFJrK81zmcVAi5LyNtYcI+iE+kn
qC3ILBFp0caRhMdYNu8dLqreYtIsutIv2LNhMLoa85pCZnr+TiEGXEUNhOvQSXTM
JWMkaY5z9f8bOo6tAr8TMtIZT+QzMN40xqRWSeHnfXJ/WoPuDLKfwmjAxXhOM6jR
kcDwFpn1onS50qn39LOg6pm15oIU3vKHn+bcFVPow5BvvdKvt57t4HP+uFKLzFja
vHRgFjnynI07Tzrxme+3YPr/U3QZv9Q0l1X7WcSAiCmmRHWAcVs5f6+q42ej8Vpx
ndMHWbT2Tqo9tnQjKdE2F1y4L6dYJOZOW0wmxmLa32jgjX6tX9iMEXKhX0B/Pf4C
dFrbHbD37zRzNwgECKDdQW8A/A3eY/5SdVj2CHxmp5o0Zbx2OUyE65KBacApvSLI
bkJFdxFs8rJvPltV3o3ajbWpHJ3CPEoW5jYsd02BOHiELyQQxY/r176UUgH/bP0z
yI8+toN+3mdI5tDurH+f63sBNWOWyr8giiS2Wu+DZAoWxOt+6p12pMQBgHpsUCO8
buTf2+glHJCdHdq00Pc7TkWLmYNgpBkan20vjLTUmeU0X8UgZdeGBtHVHg3q8RTw
rcUeT6EBYt7mKu8J34Ogx0dqdAbc0tWTbet32gnrXdlLgPfBMZtBBLvSaPuajBfT
jw4t9Rc3Japh01atfrq47TX9KUKh+hZhZb79QkAgXek1c/eIQrwZWLVzjBlf4+gT
VjlvFsvSUcJs+AhZIi1O7sAnO64aUO8yrVTjz2B/aoo3VaRoxqcq4nuVpnTJRQPw
j2uwsLLMduvy/iYMGZPL64SJeB5fkPDve4tLdQVv4+5uWZN035vZFeG4UcLi68Ux
zG2/BT7f84W8ln+VepJqS3L/kjly3pMAvEkXXvnhOZ62k8RHqOHq0t7CEtTXS0HU
Ttfff71uCbxg6Oe2rlXx1dpAoDOaSRZ/AMZ5MMfpIl6rP5/XRRgvvXYTlm0KIUiL
9UifcXyAV9g2orTjD1kDxKIqOA5cZeI7hVXQGAElJHRsFrngR38eSs7xcI6AzAoL
92fm7c0GoHF18EZ7ICGsEHWi9esEW31/lfch4P46dU9R9EDMdETcXKjDgryfITni
blTFjdSmOj8rzudd4j3XK9NDBMPTiwzryhBxHLM8zEpVCddkhDPcv7oMebBUZISE
GzD/F8sx1erFGpT3SKItBwD2qsT8+85d8MW2Ej+8KSTj76IGH+MUSVNFYvi/mS86
YoBqoIOwwYCUylHKaPSD7b4l5uDPd6RO6xZ7uNOuU1vBRXNxrCkyr3vkXlqAzyqE
618aH3gyCl/tZgJjmVsq3cK0fk4osjwEsIpIWPacDwk39xGigC8OLUdkYIYyla6+
duVG2nZEO6e4ngUrx57o6AnBYteWLRwD3202+meFbGpFHuVvop8rUQ53OTzopXOt
NIRqQRk23RXrtXG120rqeI9WuhDwktcd5NLz0PwSxC7Ivkq/w25vEwM3tHbU2dWG
hB/uFIaQ3ctu95Swcw22ttTxFIZLod7ISGRSJ9ut+0bE6zbWuiBGtnIkUTi06/kW
XbH4EEoQ2RDvQW410WTw3wpbfN3jXyu3t8dYx7zo0NW7vSKoMeDrD4ROICzzyr+x
xUhG2XWXKML0pC6HumCAJ610Zv4H7QGkhO6la1JlD5M0NOP5hF1LuFlSmmm0zjuU
XGOFNYbLD9d2aFgEmT9PT2QtmeVBm+7rKdUhun4rvLTH4AmbZB+Fyb0HpebcdAIo
QayAPVPaN3o/ktmU1Ka5jvKsarzAwAbN6Iuf5s5xS6fg3hDT+N/KUAjgrLFcrId8
r0hov5eOUpyUCysTZigJkkzH6iGfN0RVUNdrHAeyE+CpR1zmuiOHHIhm9Hui9kFk
ZBsLxCvgU6R8668kFb+wxKwuH/osN5VnGxhH+UIrzpp8STi0Le/npfVvoWMY7b9A
ZekVN5BhvqkDV8UNpj8G4iVgIoL4LuuogxwnggXo9x63mNd/3bi1c6T877zkejVy
cv8A+m96WpDDLoWcnNuLJHHZA8+DKa23iJ4O5T1KmXn0LfqM5CeggPgiwQ3x6CK6
gsQI/Een612UTm4Ub0XR/WgUABnXLfOl+YQdiDSBCYkPV4GS/Ba6MPmnn9DmBubp
ykD+Tcq49VV5zjL3QHWvgN3tth5Y45UwfKB4mnude63TkVF9819K9gvQvu46Ks1u
eNDPjkiUx7uniDgg22rs0IGGIbs9/d2grWA74BxwvnpLS7jy73ecyqxYzC3aHOIJ
IC8ty+oNbwhsmQPlSC0gUF4JYZMroFwy6PKtIa1ANFWarQkfrmJmzdmS4kLVNqhw
QcJkKrxpTCP+kn05/1kQwKwPoryvhFQ1EjJhPc546EnSydc/E3xkhFMnTpvl67tv
bXBFYD8ejAouh8jDQ3fWJ01RdW5A2AvhBdaKqqu50xbX3CInvlXw2kg76yPYTN8B
gshKAyh7gsibTwNDDGghgA6zZr06mYhYoUCsYDH2a8uahHFQsnehjSWxIc9xcZEx
J+FQhFjbB+sfUzxp+xH0Azi+7uptGg/sk2QxXYOKXNZO34GsWUaEPLj29G268tc0
2qYKjml+oRvmSxgQ9KzO4diZd7yj3sazeokd39Wvhz4HjqlSXH+zqgNchdNZ0+om
OJkbwuvrSPpwH1srZGY161YnXs1SwRxDBLfELaNfqcECiP/GojuZEF+2sFu7skBG
J+1gMj9NzbtSPB38CNiVlUfchSy2v1AfnwnqPqNdy2e+o17OQHYmYsGJ4MY7jmbW
41j3ehXqQ+vl4RWgsd05ekobN819Wm6FAaefPSM/qNlAVLfb8w57eZrqCgl8lJC/
dqu/geLnBtl/9dbFAE2De4A1YQN9OPmAmjq3FjUBPovmgvR4vlVxMllV9mF2dLa+
YICjTuVOHGfIFWUjsvTL3WQX2GIMJk2dbK3B5ByrfWkdxuy/yO+6AoePwpAIuhpj
6ARKhY4D/MTLDaD8+i39e4zCWBwPNshr8lutKYebhy5rjv8c4R2PDFNk5c6HvDjk
bYsq8i87vwZbTFXTVINYkAWkiwEwDQSVjo2AD7tbv2JTniVwmwk0ECA6Yn7MSc8x
ntk0ZAGNR1lnJR9uHFTTNZBcbQBOro57oRYI6pWMDQMLZ2df/FqOgKkAxK1rS0bA
wOBTpA4neD/nOL/sqUw+Y2qsUxgjCi9pjs4Jf9o3iG4/UkAgT3ELUe3j7utWbyLj
zWD2r/W1PXZQnarkD2Dt6liqfn62dbeQxLFMaoW374v7RbC5mmaDRzWGv1j8WAP9
W3rOJOn9Rg5FtSxojM0sksNzjzrODxCJKbHk0r55mn1MTHSu50YLlPVJmAD1g5cq
GVbcEL4zkREYdlFTIC1iYjTwDl9RWhxuhI7aD2iP67blQXcJDDgxQqJsKNqoWMHc
ixeihVtZBfY0Y8+8fXtyP4iGktG5RDgHq+HRs/AHp6HQ8jiGosRISMij+eQl/cnl
oPneoc1Ze5v2kQJceA0cE84frTRIjg8wkJN3IFsKr+doaTkzOCZNxCbfBGJordyK
F7Vkjb+FP93AgL2LhiW+UQztoZiLeqrqv8Bd1+DxrgjBQhpRmDAK6qRK9TTaKrHQ
EnGg8aTGRvHQnMjqpiK/S/VaOqUOTPQQifGi+zfxFW0ldLDlfkVcM0TLV0LwkbmL
Ix9o4jvq2AuQx9WGkrynCxVhGCYGYrpCh9/IIdysUWnk4wifV4jV6slu6JSsxDWq
7eRdwf+RU2cSMa5S82ITk94cTK+yfUn7z3oP3SmSjK6iKsvUi15VTnjiZG+IrYpW
gcoloEqsmH59Md8tBMcvFP/NqoLh0wk3/IyiDpsAZ/ejYVIRuxsbL4AJI2DVaZh8
9KifNVAJaOzsf6xdH8D3vhqEANxVPeeU556u13ouJfR+PBlQ0tlM8/P345J4gE3Y
5yhdLLSFVQa2YLUjiBhVCnVevun5ZpD1x6Gs6Zv6+4TtVKld+cpYaGU7fouCgh5e
Bhl1BR8qhekk34M+9BEw0sk8zGD13yvIraYFwrvQsfVg6KB9aP+bA8CoEnjNVKvw
0jB7rAOTroVYUfmzyvV1f4qFiMrOTbYRa+xS8I0wdDDZNlupMSH9Y5AkmrXtUUje
mNqyiC4JyEAQ6vGPUbfW3WHk1LNqjJj9Cwm1DIu96ikauc6mw0jaUycDLzxEtSdM
JuEtOP4v5oFjO+dSEwmrdAn0xRZZIZ2woWkkkGcVbwt3ZVQMhnT6qv0IhVnV4wGh
I8GR5fEHfkVLvEWbSkyEpAzopELm7y8JNR0R41R4mdbFced+69eJwXQfUS86Gl0H
cMm7AnO+OLarnPWQxDNpmjgmD07QOGDhxi6er7OJ3dcxnfT6aTPhAuZTcFFXQtJC
pstRhI+5WtAJjQn5hiIij0C7TQpZU7ntSPXYXLmh5JN9SsuA2PRU4R46kM6IaYj/
HOcquuWHajG1utxSNmMoi6jwlKcfz/SS9GmkROo19ibQbR8chP6Qoikg7m4M1cN0
1i9Fqd14ew4Z7Tp/uDL3sfjgvIm/srioOmZAJNyEp2sMXVnAhfdbybdv2xPnwTr0
Ml8Yat7ChK+CvBpnCAdfK5xb+ZOBxUnjBnu5NFNRuZuLu8EYnnBSPAK0Nd/73bfK
ktkQJdmuNNLXhTluGBzwEgeYTgW5jiCjL8BlTycR00IhmUzxyv9KBjPKRPDBVKjg
2+fthXB9XwP5lGeqxr7HF/HNN2szAcJ763G8iL5oaiC8aNgeIMiMw0ZxFc6A3vD3
ypY0KPzM/GonJAHLBshDs8fcIqq3FrBJ4Zkf4iCL3IJ67YKCcCxaZu3Nox8EYtBZ
eew2Chf0BBQnssLFYl/q+38v1RGTbg3c0WHMRnBWOUo3BMUuoWRfl8tDf3JcGj9g
uWhTvc6XnWsU8MOytuY2HcbFevtHE/AwmQIxFmC9krmZgPJpxc09aUMv/03Ulp2a
EFyInnpNHGSntc2zXSgOM3s2x+edyPK7CKzDS47Ex/J4INXEoedl1Q9s3MdqLjZ9
v5rObxit0Wy4EM2j6wrjp3DdUaQhb6sFiLfcVibndLrjmIC+mE+NgYRlEh80CK6D
x1XLy0CNjh31r59wO9FBT+3IhREC2JiW+xOpLsZ4LDLUVn0Gor/MDy2rxSUIdx7w
50Eeq3z3Tlud8CQs5nJ+ZIVoX8me/47wvz4RAurmURVpKK1iFAztc72ZUdLc1DUv
q26Ua66ieQgtnmSa2OmXhq6j2IvYd5kt+hZOmSNbT5Xkn6plgzJ3aheZuq/t201C
Q2eCU4Calbvqb64sAejKPi6tkblovG3ofaaFA/tVbWc++KD0gS6fzr/7Q/8JzgNQ
wYcIjobbaiK0veVbLHx6L4ZopvItQlO41dqK2zoFOWAgUjmPO3H60jtgjtgK/lfN
4iMB2InlGRNgLBQiaBr/IHOuIeGu6o4AQq+njdJNS9fop84t77muS1sLahJ9Vnd3
VY8YIwXiWKKT6BfgxXO8ENRPLT+2zDchfiQPpzEoOBJrNscvWDhqXFWjxD9ZHpRc
edcHmi1XlSVM5sSngirAYJoFHdyy2t2dVWf4W6PjcUFoo/n1AnzBUrwbibMN/cLQ
jhG3H0JaiTc8AXwn46ECBOOZMZJrSSG5mh5oZFNxSj3WEtrBKy1xJYaeRjafLrRJ
3DjuTQr3rj9hVmFmN7/HUL24lAkpgCB41vWJcbfAIFpqEAc/zCTIJQcQqvHVR7ms
AfSpMc2LkfWD/7GgGsWktUgb3q8Z/wtL+NkuETGJNdFnvLAlnY/i5TDLvttyL/XU
vHTdzZgxdaxZCSDFn+pR8h0FRBmDp7fFiTpNw5bLoLjtfZ69On85kGHMUg+JFKhv
jBzwGV8oiRx3CElyIft3oWEf9LuoVnRp/Xi4gwHDj2hkwrYcJ5qz+eLALBAJNGL5
mKaQHhUcgs3xQTFTFC3hbY/vKqI7rE1qLiLytVd2qN0fDCeBNgAlXHWBRqKgdJ8p
/LZAmm0Jz/kIfhCzL23RtpLewVf14/vSNByF/fGV2guW0gGTtIUxzwnEXIX01KoQ
XfmpwDG7BKum1o7ZX7fmZqGwoYrkRTRYBv7NBsS+m9xruLI4cVY+7j9cDLRaSrix
wIodWWo7kpAUnDeFuGHrVj8oDH5R3zxSmXCYuO7fvARMkRIXQMeI3LhAtSRoySms
KVvKzTyQhILiwZctjlCcTfmIkPvgr0L6JEXhyo1pG4CUaLptvC+7wRgD58mOzD+n
/jGolH6anHfe0kb8foFeJ/QiSBdP7V+HBmWBOMF2jTn9QHYm/TQz5V4Ucd4bJyOw
bapPhkRlbBM8l+rlH3MJs0wrXGMa4CdoShA0cWsi6CbILJqqSO+GAfGztLwU1PPc
l2rq0agV/GQ4llvqUIKofGkKkJgZhUVFQ0fElHn3DfpBWYl04hYEefSzyElEcGg4
Ww/vd3BT7Qeg1Xi0oPLuxnOaORAKl0tfMIo0YTiAED6qEgo76n/M1JJEzIJpBBBj
9wquWyYxReYiJccPY0mIGYgyu7cGR9dCw/21GMwfIk+s5kwcaFhvdmImGYNZe+oC
JO05vCGPSmT61KquWgUgI6VW9tTLpxtzTRysMw7w9Ke+e3X0tH8Vd1tbOz383POj
i3+s8iETEcDM90SzcHcJr07zS4EN5iZjcXIv4fedccF/a9EnnCWjC+F6vmEeZ4Be
2MczLyUxcQgfpLikZVj4Hp97X9N75Q0Drl7ofvQYQ7Rp8Fg8miEt4H0mNW9Lwdo9
qt0yRaBU+vVUzkPnVEJxBAUzRvysCBR4RKeXo2xtavUsO2c2DiXizOEJYi2jrvQV
+Y9elZLc452oGQJPTwXUbKwxyFvCpe+fLWRdSmcPPkZr/RkKihSiUtqLJECjdIkv
tWM75PPECbGxZluPVtQz/mmG73cYavc33jutw/xpnxk8zNpXmb7Ij07ebeqMapKM
ky7SKbNUPt1fO7ywo521DTMjH9GIag5QmNPgem9CScrvwnHm3ZYwb3W/EplujdrP
veIcpGmhGKsroNITyFaFGsMgMe1Nw0p4SXZqd9OKwAN9vWvzy3Kf6wXgvkTZyTqy
BwV/syYZviLM+ODEfJSykEG9oS+VcCBYtRqGvRRCfdpDT378ZwA5pZEtkC9FjWWj
nE1lbdsHzxOVpdNFxSEwsXXy8yHhIJVixt2rOKGuPGTWxAI1qTUx6sAgVEjzogYd
r4cEhP+ihWXNBIRvWVIAxEixLYsmG3PI64ByIYr6dT5jrmYfpJ/i2IudgdS8m2lQ
E+q/ekpbyCEyGJL+HSBvJTD0bBa/d8rqzP2esJX9uQFdbf069NwsLVUHHJAK8gY3
HcLW0Ukn7AZmnhQYiUgacgpFZViNqA/rZPdxVMDXvHHXwOFojABqmSQEYqOpBsEA
XeEkUA4EJDlzN8p8WibkzBiL2gLSSkP9GKrBYkF53d3FtLYEzNHV1lPDjCvexeZw
cZcKeJuL2e8yqVdCIl3/ME5p0WPkb98Aq1LO2rWMqYpu8WaE/a8fWyeqaRXbKMXl
8c0ggp1R4OEDLnvx50HOfhZr97y9ZihpoldYqg+qLQtKRV4vcO/pS71q/NmXpXA1
Oo6sSaw0nVWJgWSxj1H1IfSd7xdr0fTjR4nwjz2+RQjC7ft2v5NFqcchyaJvqSQg
wI0U34dcKseR4lWLS7h8+mKtcPFp6XTuIWzds8ehJ4KPwtpVXcL8rFN11CAcvUiA
183ioIWSBIXI8rrG1W1bZVLtU3CLt/ZpiRlMh25g5mpqNYKk3WFKgCWD+iJ5KIK2
D8zyWVVBnQRpxqeoHjHqVAH7W0LQS7rqWwh6RnsotuFWBdzUbAIOPwrYoO4sy2tl
CUIYk9lJPriD9GdAVbLEAnOyk17QOTnNTSWe/JBHdpPnZG4+EFOgjZPC342ogX76
XL5EzwdYKiHkPgFM9kYGixMWGF4HSl5wOpE3pgMmDR1a89ATCZzsSgvvgt6Z1ob5
TTo1Rw+OajtTYGZzZeG3Pg95MZ2qRUK6Tlb77ozeQXQIjaI8dkyceMFi0KAv7NfQ
AbM/t4r4KkjbWhXtxMV6OE5owZ7FDsbm46pj41gSVjYjUsvSoFGgsS1Oy+nId85E
RX8B2QaHiYfznUdcif3iMdb7u0FYJsbHKzg/+/w+NrT3D1ZTJwbEuW07+4cuvAbn
u72ge++vqO9VLEksQ+ry/G7v5gYkI1vYssGX5Fp1MvnwkZmnZ5uy/sOeUvpTnHGi
2ygECEIkkxtDKN1QBNl2hswur8Ei5Y0meHmSbdudW3seqJMTr8h08lEycw77M5Ay
HW/gvmvqmwCTPhJ7sHkbcC0289BnhgUIuXzBz7R0Cg0k4HNZhekGPwfOJNF1Llcz
PSH+92vqCo4I/9puWbokfMnu1CoM3uyQsZjYJ4lK7ko8sJglfVykdM9M/eXOCtSg
qm6Poc8oy6/VsIMiZbkKtbEAbfP8S/Uu5gXJA/jW+cZpWfu5YQ+gCV+7FxN8+xKs
KTJWI56/TdtrUbXsppdSAZ085SYKvQvzkkooaJLHZC5RyWmR82vqEmFr8iAr2Mea
O8xEPWYEAkGQBWv4rqyohgUcJQyKwvodYn7W3Zn/ej3/zf35vjG/ltB1ICmNhyRF
CIdGMuxDla6SyRtqtDRSSKPgUIBsi/CAFLjuARB+RhzhAmkdZiAQLxhfA0FIfUE6
9elWq6K7QERZdvwFs9s8Ew6iQuZNr96jQ1MFFHHd3nHG1GYnESTbM5yCJG2WZQds
zaWvNldp3a784PyPGTnxoiq5RhL8AoY6g6MYkHfnEjSOylmBpkra0AxiWCZ2oN9H
PeWjbXbpKoWBwSUMvf4/GUV75TXzMKE8GynIPhDvYkHsqxxfSmp8h4kJT7B2b42r
q7HRclogWWMZReQQkH18z+Ew5E30czDUypLjMS0x83Paz7Z/kAsZaZRDnNN41KF1
RffALBvmdE4+XMi9x/t94IO6Xq9YOS3iCteTAPJJ+sKg5FHVvIRO43qspX8Dmdmy
cyIbgYnBKq88wY2iGs+4fnfhFBWSeG94tCDNEaIYaOPjcmN7lUCczfWbwMfFwYRk
qey1BhtzyMDuVvK25/9pDuj+pOojzlcIrVo/zTd7FwuMWgFWAywNOANpwqtOIYbw
O8uSr5b5nPJjW6cNDoJ7FqNPyZDzC7hS4Sdu9HUz8wJC3AVuC5TcTiiFVYCb0QaW
dbAHF5LJ3cTOI0f+EU8OsTwMDhtyOHL3GFvyzi4UBnnkWXhPywqIEkLT96lZe/xR
6kTiXJ1f3JZlE6mwGFU5yW7hc+0SvIa0ugUjuUMGseIkhBWqI+Kq2K9Gq+845q7u
H/vGpDiaXdcUEnvnR9AH0TS2Ohk0n6Q2+Z1d7Ukfx/wu486EnY86T8ekpGT0hmrl
Wka3wZsgLnTpno3twPdmN0trLB4NlD3C4bG2g3qYBUGPdVwrROiR8+O9jG3Hmd2v
ZE5p6Xj6bR1pqYmMoMwvNMkR0DjW8X8gjexvCbmJ5AL+zbxPM9aMcq5GpnWoDJAa
Al2uA9mUcJNkZ72Bolwby7QLCImI0UPJMiB0aTyJhMbFIIjixcUf1hY/I2Vll0+7
QzOgF9dKkDRgQzeKCKyRzFFCpLG3tnwPTvdxYu/bI3aNyfMHwHbgl/DN4LX2jlT1
kjlJjTWSZSWEHf2GL3byJRuNQJfe8q2YXEe2ulEvue/NJ0PFVrUpV2SdTp3LIt0Y
s0xjRKvk4STOvJw+cGm/Df6ZngpmZfYOe2qieXEHvbs1eVbH8EKO69fURtIyiQyZ
PJ3nSNItdzBDesJTpDiVKjkzMwGR4+vw4FfUwZtoCw522zYPyZwRCBTdTRpnbNw2
t81JrHGpI2wyrlXZBXOICYzTGblvp4sfnrysLY+yJSK0X7YSPhkaBg+2TQoAkL1I
fAcWBJMevRbtMQ9E0B47h8JjS4WVlEN7SR6VyBCCYLsbqM0VsjXkiMKrAN855GC4
4rSE5BGrSrdcpldJABSPcn2HoTYlaBR5IbuArgURBD/qb8+GUu2kWzgvFCiKTvsV
h9drPU9SGMN6jTOB8g5hozsb646rj2lOUObkqkxqozT6o44dKUY7oUbqSbJKMevI
BANKKNSM75K9AwEQN993W6U+t7Dx7XKgvl4s7f8AyjLakxyZlPio4a5ZgWnnryDu
A04BS4fDFk4CW/TUw2+x+uupf11KmiR9IHqyhgBrC6Mls3jdj3v8vIwkKAFOO0ff
YHirxpC4FHnb9ZZOyTXk0XU3K1+iROAtu1gl/QG9csj6XAsrGdgKqnrIOymFJ/LY
/AzNDwuPEYrpNJQ8yt/hKEnmn+gVbLUxkRsMk9AiZYtK44UVf9bUBMT5ckA3RYyH
LHsZOKq+4VJcdhIGKY6en4cXjIql/L0tVM9WgyI4OraYJGsHC1oT9XCS+nMYq+0Q
qpRZKMR2GF4BuCxjU7TPzMlAAegseF0J9z9VExaF1coV0Xfv/hW9RXNzSjUWuV8I
BuW7BkHojeegG/Z9qk5Qfew5R1kqVTMY92Q767oGXUKJ8yBrffr87bCxixL97rNb
49LECF9cu4rcPrVHN0psUnqSH9ZksPI8xAIZQZwAK/YVaiRP3P2Ga2vsfRuuWB+p
Ua72cgFPWdZcl2V5jU/+IK3rwSwk3zOxvbfZwKdjkw8ZHVsaBz7kzUpeGvJAI3t5
oEYT/jZv4lP6selUi7clFao+PO6fWYDcmGE9pXX6o2BaTVoDCtFj85t3YvpqeS4O
P7heP9+4KLrZ2oxAzFVX0hNUFSnliHdQB4GXEIBINfu4URVx3rAZKsdxbVqV4AFA
+w2gyUX+J/bXR9uzjWIrj5m24MT1qrwSMSZtR7vA6p+Nk0s+tQ8Kwq1iq8VoCQzp
ZHqAkdYq6nsmf1U86IWLxUHrqjzLKY0A6OKMw33vHY0ZRONba82lOgheZoaiWTwV
Fw4STHv0P4rEboKEkX4aJPRHK/Tczq82qAuICYVkaL11YZD1GurJVpEBUa0y5qLV
gdFEG/f0P/CW6Hr2mPP86DGsBIwir2Z8ub7/sy6t3sDgmMqN8nEnAhIJJd4S1Uuz
xVs3gka/118a6+pTZXQVC3N5ZsL6jXL09nPa0+BpTSHTJEVL0wqxrondxnudhLzJ
4agNudfHA/0akRmlrFohDIuOrp1PZjxKBB+awguz+pyareb7e62DMqJfEbk1vUQf
gUWZtHg/5ufcDDtJr0jxC5kFfyiKWT8prTRniTWwiBihORhfzeQBKFH20cGzKrDh
l5tneswKc6EWDoxNwDN2TSsTEsUh6wxrVmsnYPlXTl+wTkGzgo+Y98VV8pz27jFa
9hNAa1uXdPMeSOjRjSKOKTLhgE4f6IlqxJbJRfEb9Jml2nM8YNkT0c/LBulKu9ym
Qo6zkfbtQ0zKYeXFbcYIcYnaeiY18Iw1X+OLUuvHiAAgYIDdTN83lsJKGt/4n5ms
2n83ZVdQVGXIelGJc6whD55p8hJ5rGJY6kkTM9VYCmrH8FiZwo5lSRIMmSja2/UV
7lOWlSzpwroDvBHQU0kPBbKYMK07ZkmaJVBesLIPI8FmRGQzBnffZzq4uELAOGZO
md6JDKaLEFPdvGzYpm1P1fsdGEdAb/Hs0tLuSHIpdNfG1qJ72Q7+rLuY2Go++x73
cnbwDtuaUCm/rF7N9GWVRy1/QelMHNqWT+fbCP/GmV2eU3ZlBcMNpYr2ZFvZNuD8
UhPeqcT2v3e+dGHHlnxqCLSfNw0NwI3ETGPO8IyDsY/gmE/EmoHyx0QJvyNX0VO2
AQld/9WwCKh4katu9CD70lcYOxnav7jKDdNy/sRH1vq53vVSOYEA+Mc33/cgvIW2
pHnhwvkkeDL15FDsIGUeiTBi7sgdvveDHs2pcA/Kehl/PKh2x18ky+q1D7SFK9qd
hhRhwEy+IwV15/kZb1aHhbTPsV7IdZhHXaAlGkqZQevSzXwuX/NMOqLg1Sl2+3+4
ARO/zgBXEjblgMVxqh93q3I6xwd4KQTWTosYU3bHUO3cz+3n2vUqonZq3H1z+sF/
46eoFENlx3Mf6URD3wS0MLZMCxzSIUAXQdj01RoZKieBGWgMd1TZNMXCnlLUmXDC
NOQgRCIojv6DP3AJjwOWb70zPudtxF6s3GxDxpEooh7+MaO3Nc+xsANHbPVAlZUF
KTuZZvyETWIiCjgAxCHyQiVhAf+5J/6p6M3Fcm66VvrTr9aoZ2pGe3oypGS5dQt5
voXCNKJOJwIq+kQDjXpdLKY+ffbs83R8tPfGtC6MDo0nQASUKw6aaCMDV1DvOcuM
RH8nqBtNo8ZAPZuTaj/nlaALjNlN8pIwBb2gt1R7Bb+/94ALPAiV1E1Q4phwJb2e
dIqeP11tedg8Mu/umy/y26VN46AQ6BbiVD6VQU7Ab3k9AbhrVA0tTCsILsVB7MSH
v5EuL9PjaRDy0gdUpG3uyujmDoQ3InpumuKIKSiYG5AzRnMH4q8s32W3jR7GfvEB
yNeUeHNnqywMZq6/XWwJpG/IwPBZzzTXxiC412RKUSDMFe3EOxg32xRCzEK6I4Im
nIgrHGNgyq/+Wz7YuyXUfWchPj9M/wMVUnnwS9afVYU9I3YZLqvkc0NVLE5epO/t
D0nxT9C3yawV3dkwWxEq5aSa7JUar1aWviuxn3hJf5pdyV49QkA6kEmuuBpQzeAL
bE/MxXwK0arq8JviEBPLCT67Kr7gEyZKo9vdQZ1RlHn7ndQ4X4Fukk9qNM2rH4rJ
cbntsY2/Cf1iM75m7meS+QCUiyh1RdZsVtye/5tBtpwkfgExFrWOH+KEvwxl0PFn
ezFDw7aQW41Gm4jy4i5xzGRa/3PgpeSA6Vq27SNqcwP7JRP8SGS+aJLFQyqp1L5H
OjljvrrQ9K/TPfQno6cODxkQJxDHiRtslAHVvLX+uVz8Jdu+nbVy/jLjwGo/aRE5
bQqtBYPHoRw/czU961mICbXoU6Ke0w/Dba39ZBC1W5+JkuXC0JT4J9Esh/r49yMO
799C3ez5SWhSWE4pSbRhRgXDF0iVdZ54ChEFvAkqjtvXt2TQEP143aC5BNWXlReC
z7qk7VhwWQAdVlj1ZQKGbZ+pCINHcYmm6HRJv4QGVu06qgPfHKifTjZNWLp9PDuC
I5W/7TQIOZlAOdV43yCxROykoOQYiRCsfyk74K9/KDFTG9g3/Qojp7kXhe/6iOCW
heYwf+ZECnRN1We0TYQH85vFuIWbQpWvv5oQ/uHgqQyOzuTrORlr407ffQ8JRHX7
WQ/2uJZRe47EQpZE7auS3YLwcz4irKV92M3eLc0QDeThlJCoqip5poaXV1ayGogC
sITqJmcs+yXGwH6/C3Qek5czC2jwrbqCi/YDEU+j3KaoV00IrjoFBPq3tz43lf6m
tdmN4sMd6UX53cImR6hK4rmiCqiHsed3PaeuBXa1ekU7bdSzMByHVrRxtS/p4t4p
qD0xQLb2rPOTU20Gp5qjTkPAICu9anZg9d7qGhUaa4Z8D/ffDcrxWwBywR0celkh
shKQb63PN3o+64gb2DZ3trYeIJDljCjo3hzs3USF/wGtQcZUpTNkyJyCXxBfveK0
FLLk+2dHCD5dNEVZl0bhMtoc519YVCiP5leAXYfFfAfmv/MO2Lr5P1ROpmmsrS5L
R03omeWNpE4qVg9GvoDRrJkp+V67cP5pKtD2ObU7YOL4zm4fRHwX7lGkCDxN1GI6
LZnQJGwjHBn/mh+0J057hMIra7AMbO4gar/NHIEsYUT4ItP32aveurhWAbPCJOMt
7PYmrv5fSltDO4cunSVzwiWnrHA/EzxQ/SHCGTWlm6l0rNTlzqPEnjZy9ekkO+Fc
ForcKuI3pPgOix8EZgha+h3rScP5Ch7uGJe3O/bDidtVqIlxx3t8dA4TP6OVZ+/u
fMW3zZzm0cu0TTPyVzYiZKSA+KwG606KawGep9m0JJV9EanuHdWhLvvTd1kJBzLo
XOxM3wk3i2BIHsuAvwEOvsCNWesNrQjmzbGPEl0vowhoCdmD1mJhui6itCvjLpU4
HkhhD8hebaztQMDvzwJrehGVOo2MjGDGLyYPNATbnBJzbhFubsamT0lZUS31vzWI
GxPo8cFIB8VMSn8KwjHb7SOl+5EOgoo+gNFPwewT3Gi2LJOonEFT8mpBEuqVSguH
DPaVbpxL1qIIuRTS71F70s1uNXqqRTG0MnGk+iEEm9T0hdkJnDTA1VQ0DzDMbhTU
hUqO6SZXfcJGr8I+o+iKrCxFDVnQc1TUIiyqdG0KgVyRmnbvnVyI/o5p5ofTbYSf
ml87TjFrRzR1udS9M/zeoDHjnskbg4EBDcyS7sjYz0P9a3brQN/6LS3Cjzg3w00B
T8xLNeJOfrMdIHaqiGMsUSL/qYEgSryZze71pwMnyre5GtnSzYphDgEzoyb3ZdoN
r7b5SWZBWRtew/VpXhsrTuOefMzYqwctFPEdIo57EzmpPiheMUFOKf0P93WaJUKv
Mw92/SbP1yTqtdfxByTpLnSWdQ6F+oJYFFdN0Wi+CBQ4Rgp+jVeD9SYbyOEPT5v0
dtR3BNfXfKM5O1wimx7NcJP7NLP5MuXrCAengk1c+Ols5Vc6Qu8dOtCmd5LtXBSi
7MvqigSDVGw5F57KuDMMPF3OvVTOnfJvspxP6YrUhLkScVJOeCEdCvBA+hlyoMPw
DbMhlVCqTYENU40pgB9VUdXZ7ykXUDjVg0ySPFi/eLKZRJuGZrzcXVtc9QbCTk3I
3+fCo7D8WwtOfokCkPMUNz1M6SIPazCMJ9jPvwxXwzoqKkT/k2wUAs/m1qnFu3Ui
tipPb7YtLYbfLcozmT8vq16eaEsIjQ5wTywWaZukdSmsDjUQO/f0BpmzdDrILq6N
Yz6JiotKieMguGLE769WhA==
`pragma protect end_protected
