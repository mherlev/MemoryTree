// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
W8CmVXQfAmNiekImStsgSEKWIROMCvr5LmQ0LrPM+1vDVJUDr+zOkqiu6BRpP0U2zq645C9GalZX
PbTl/3cgGsMUGsGLm6jS/N9al/0UpEltrkK2a3vkh0BbbiABtnWu0wlbfjvygsvxY3iqb/q2BiuJ
3XdJ4BXTGQ7xSi7/kogMwNnE67aFYl5HJmH9AY+n827Gahha6NG2ZikLa5sRFWD+td1pCtxJM1t2
/eDE51iDiCZTcqOix4d3BBiP0ioi6ElVMVrb8dhDbunqeWsHmTqU6XQepeQ51w7+TQrVe1/Eav/O
yiDjWZHbnjh02sUDHJdR4NLr2mepcP9oGMzfyw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
Cget/gmKX0+/pG3ZvdUPof0IZp/KAj/wces9EylPo/L1PHd/F1KqEd+ONDinrkCkU4GGohhvbnM+
e0gyfqCk09nl+AIGzX+7xJuvwCoDfIU63yte2pKG6yFZQu0jDEHOe0dPxprx5qCRXsOVGGy4aETJ
ooWvdzl8fd+zR0lywvR7jfTENzYTLfsCwhED0ZAnzrxF4kBGPyBbHNreDSCfWq13E+24xWY5cdmW
MN/tme23/yCd8OYnpMnk/Mqcz4imk0vCnpo3ldWP133TSyjpvqGSuacuN9HUJPNxoCWdEyxNZ5Ok
kP3HqzP365bZipMUIa4qJ6lPEcyyDSt/nBSVbcF57hsxJGxzn4Cg140H+puaP0AVHCH1dFE12aPm
1H1ra5y0sFRX1dmov2Qeegi6Xb5apgICsBmyRqcoa+29omhRSt8peT2qiJOTNn9D6nh4/gZ+b44h
r3v2qsnDs/NUylPP0aTrrYGhE8nCgx5mjlO7xO4xzypVQj12/6UNGVy0knb0m4jXweaBj8Y45cn/
csL8Xdk1OH41vinms2jrOSOXePBsMebRp/SaEMt/ztFT8dp3o2z4fxLym2sSbcDqUFV8CBxejjj6
HQg8n8Vqu8RnQuVhm9vYQyqYdwBAnmWWM8sP2Ou1Vt43LRjTKOvCIncMuxizPR61xqilIJ/HZjk/
I+IkGSpTS1XcAt6ERcdK3X5iVSVzaZZBvEZ/TYkFCZEIxLbc309qGWhHOh0GNAYnKCqQ3EJH8EdP
pj1quEKqg/RD8jfmABkyyvN8nNMcXL02Vefo/YyY0zXCZMxhire3SgWrV+fo87UPgIMFpf5HxZ0Y
SSE2fFR0sI4nLXZEAeJxWNbWt56Cw7cHoyuyK0UVelyBuvNnvIEi40XhLJ1Cd5TiIyujI0QVFOCo
FMYTSt+RnV+01VBOfcPDsiUH7f78w0RH1DqVD89zBLqPFhgVlhq+7sP5VpLgBCa3H5udl3UfcgMi
TBfLxj2wku0Vc9V7PsO/c0hFQBhz1w0CShyVbXLolQMmMM4xB/yazdvKwsEQm75iC+nBKSdn2+v2
tKileJMSLQ2uuevLVUpXCvSXgajP5MnjUzwWCR801XBNd/BWc9UAaQSy4vjcSgD6XSIOR7Z8gaSM
eee0Vk0WWFhzMIpr/XLxnZDT2whK4I11oQI/XGI1LxiKLUAdpuyB3Tw5Txd7jgS8eKnWty8S8nZA
T83zHesWJYs1cHm9OX9YFEK+ew0pa2rudF0dyBEgCbvbrcYCTOjIN4Gu6mJAii6WOqvGA1e0dWwA
sUf6770GiKJhTiR0NnOyYLeQcMwK9/kmctDdDpvoAqMEgOrMBadKcB32BRPZwwKr3VQx3DdjJp3s
anTXdXFbkcjpbygwA0TMdwMYkvyy7R4CWLZX4UnDxLGFIVSt8hmAr0CrHgf4IE9iVv077g7kdE/q
6nYDXT/auhD0s6KBZC/WrRIdq9R2i6qR7MAH7TZ/B2At0Q0XDFGjGr+arq6wDRUtLORs+EjUp/DW
NNB/oTc1Garfm5HUNMOzDvhUIjeP9wj+FJGrAnB/LVicoCFQaqvQe2Hnv/X3Z3cVp/surFXYUeGv
eTBMA8A1WqS9GhtRPwheUXl/8fOLwZ82628MKO5ZK4cYGz+SPEiLcVk/7T8DfIK1tUboN3wP+x6R
FZi/Wnf30wkOwm2FLEI7/PnFAg2BUZ7p0xwTlU/PeM+OVYQnw6L4czu4L+jBwZbhjkv590lhLeGk
wktjJUKk9qFf6q9PZpWiJiVNc2i2Fi/TdfqXQxE2WDa3WMPjBxqVZLipQX87vLsTeEr6Yf4fZ+bY
lQPEQa8IDBH9+6njS04ALV/aA1dQr6KoouaGS/ai8NV5a3yOmMkwJ5D1Ju/ShxYvM+SsaKWpZU6x
+XViNJA1tvXrrZrSvYCRB0jmQ/cP20tuDmMkcgthvGR9FPO4Ae1oILRCSuhhFqRdO9nqBqrIC9R4
erY4/cXveVMmCg+jcpdBRChp9MFRkS1BW5saWauahS/X+ySMs+0YofP9LZaUHv0smUcE377WTvJY
KO5H1oye11SHiYfdNDhJm6DE6cWIlr80kglcdAn/dtoyd9+iQEL4HfYK5nSiOx1+BYX41BtdAlF3
xGjQwx7tMZVWnClJKza0c93h/dD06o68jGk+WAFmTt8mJR6hnjsYOeTNGq01WCFihntZAy65zo02
adIBeQJPu3eiTUu4KkeSbOep4YjEiSGaNzPeuxnIbDdPx1dIIYvYDs1iqzRb9fl6JSVwM1oat+9t
RUdR6i0qGJuIZaLHUPQL1eRz20R/EsWpfyLG4Nn7BOExATFVcYdSQgVFKz023zAGQeAqUuZsNVtp
HaSk3ERY9iXN2OvPHv3K5LXQbCD+RqqT7elNb/Og7mcQVMix4znRigOhmJQGQXFYiaAxJxjz53x/
RknLUCW2paCaqkW0REKaTQcOTjfxa9U6AexxY/na51jzzH5pgMRgABNUXNhtnFfXqDr/r7icDsaP
mEgAkhKtG/Ajs0ELps1leKe82fiav1OPS2vLYiPKLj/IBTQCxIO0ZIduv7xSYSBwkkpwVg6qtMIt
jN+cbXYtA7mtAmXoFYz6cPqMTY/E0Ahpr9YevTkZQY/pACRLy+HtnkNR63T1wqiR80WATzfsnvY0
DZneJY9yD3EjkWwjqMiPJ+bF7oyTZBAG//OgoM/X4SWznIrNIUmRTdPW7URoBl7eicrWZkQd2a9p
nnLnAUE4UyRzrprr7XUCkVvRGdpaW9EtMn5YVtfxlptsbDoSG/mkFqfNB4x0etAjrGO2rPV7nV4L
Zw/A363DJ7gUpUxHOpU8/izCG1mLzRhErNpvXzvLK5YDk01e6yrByRQ/wjQB9N2YCwyfBR5ni1gC
w0x1gykN/sEpTEa8PLCs0IZ1CrD5lPsn7LVxVQUO1jUh2xFTE4ScDw5oeJOIK1Dp71i604dXDMEX
ZeWU1hV5wtWiS2f1LqWsXDBv4WjTgW2lXBV41zlvobcVgHHO3xZszMXnDUYxbzurNoQlXYb+nbiQ
15hThjzUGe620cPgwOpwBqNJBFftHiqBrEH9MS8v31ruWcjzt2Vl9QI0WWWrCkzY29OIq5ybUfCm
9S7HuohfsM7TygmJBTNTSZTc4KO0ehZW1CN2mz88MAmBLq44cUdsmkQbv8mtYptfp4Voxv8XwR43
bD8bfjjbT3eM8NkObL4MZpxrfPkJ/wARpSFV9MmzUzM9FdDqXkwlTCv1ObLHBZdN4i/BpHH31geL
RDPP3YiKdM80+aSnqB5eYBJbeh/BJq7KUsr4QtMvmUS9/wOBQR4yhzYlkxnCRskzzTSLFDJgNgQX
rzEiPNOOJmNG9d3JbOMl8+SCdqyCoCC9w/KW2xgJgeYtESgBIaGCHEaHSDxFexb+DGtGwumlnNWj
F4krP3GVT24hHypWWmNP9eO945Xd5sNfD99+YgtoFnzy6ilHnWKmQL68bYh/bIzqqiMBjN6/ayiJ
3eWRuXsmqIu6ozX3PfQWCbdtQgWpOgWLdmZzlcPT5rRsSjB/yJJzSEyudgzpQZ247t1lMCzaUw00
EUW/7/xI8Lp5XfHFXg05qoYesiEZSnTA68F1ZqU9kGCV10w5WFpsL7uIdoep5mY+Mgcz/Bk8Wpjl
mqIN0aZJOg8vz84PORbCn4txkH7bWRdIc9nM729kROk9J8a3uXUHaYv73mavXfozZwP3vCgT/nhI
wL5vD0XZbecaRYTP4nhScOAQx9vUVggkyoca0bcx9kwgQMRgpSc0M5MnEcW3xpDXwTDQVXopToll
vDNtFMWLP3uHxEdnYQegZXgO2fUEuE1maPQ+zuOUdFRlwGEoa6ULY7mGnUcBiCT6LK9Eey4oCjpY
uCfJ5ZbQasVM3sdP+rT/asMDHF3Yov7s9TWljh8J+RB+NVZlKpyWuhA4ZCnIeETWBrfSpGHyXJQe
dqnLJEjWCTgzcoG0Rp80TLfvhxkJl/kT4mrWmNLqPLv4AwXzcaSRXRNdAdlL7XwTV+AYQlQgA2S2
PJjfs8oSb/gNW/wUX9Ln/IoTbsEx1wlyYO3lGe25VTWz7+tZlknCeiuTRJ82f3fxqFS0bngpjMag
Zo7vSgIAsJsgxJvWOjoI6xIcPPN1oKZqahH00KGLzqRpp7z1TP6Q+midpc98AP5a+oBsHN2o5zBr
7qoTvbGyyzD20gNkQNUP6K8RqPkgrzR2CO2s+Jz7BF3C7R4rVbsiFtPWb1u7f7b35zQ3X9zekgox
mY83eoRm+SACUCVMsr6QXKbkflmnMGPjeb7oEXrEygVkywtDNb2rC0gfUw6aw6ZhSsE6hiFTTTEF
M259JXsdYQEswmY7zmaAMf+waA/NJJBaPXR0hhGqfDUjpJfEvVhHK1wa6/Hs/FYg7YVlHptYMWZf
ev7+IfcWYCQ6052nrIprVUzbOfMRAt2vh5zyQjJUcIlNfNoD8ycOpXseW/U5rxVKVvsDdq7vAYOI
fAtGahYBU8/Y3rtY117p7+KJSyFTYLPNed0BvXTAViZ15x+7njtaeQ1rtUAmupGraqIOiF3jdJso
mry1ZdVTe4vMZ/bK7eeYTYDpz7H/PhNZY/SPy6eplUiHe0aatI39YOQNsTNFMWfvvgoaQR56umED
ZiKwFrs+OzTuAkRxE50amIVXbCd9IiHA57bmGJDZB6GA65+lDLTJrcwSTUp8JnJJeGKVWk+Jfa50
QVhPK0Pfq+8Ax8EL7JAsokqhCse55TZLFtMr10rmFLU3KFN4CyjeZxstO30B8PzVVLrONdwtZAyr
1yLJSLkblQQ0VZGKkY6geb2nfvx1tWsEbAlEnCzkv5bSucgR9NKpPOt2bsb5OCEifTAWnHU6Atza
imDoanvYQTTWMmyV4FHhPcwgcZ2VwyUJ94r6R4xGVYCgplpof58ydDEF5vCLGGu+otto0ksMWEs/
sMsxi01sU23lfmrOVfpz2ecap2gRD2tx9VtNXle3/45rRihpw2MbZCnGVL8A7mPG1xVoaoRapqA0
43VXh8w7siS1lupzxhgpLG7sPUQZ+/veT5Wu6A+W3zgSmQNtn0W/MaXgXfz+GPWE84VFB06NP7+B
acYFcbzoFxcNOdVcPLw/V/UBzeqSqTrw9Xvo2v6oxicOY04GRqcWsV22iszD8U2evGiSGgFwv3al
nWnAa2VBN5aSRN/eKCOzl/tdbOz4d60p/stnmuDs5qA6PKUPlWsK2JZdF6ajTCGPkty9L7AkkoRP
upqUPYBMI30L5/fvb+9AF7E6wwc/ydASE5pLAZg2jNRvwVBT0avfs37menidfOG1AQBecueBQr9y
PrKbEFSvTSU9Eu5qNgq7ZDZwt6K/BIZR9FS5aphtsEZJLM/1cxQ6+97FCf9jZUafjrVnq4T220I8
wrBKd7lJZirpWVvododjIlZgyM5fjx821NqRqI0boBueSrdDM9d8+Wo4lMrg4cRPjqIi69Mu9jfj
Zq+3fjQ/2jq1TFcogEW0H6VUO9G2RFMDByJQNwQXp9DDKTfZCL+ZXL5WE6q2Ymo0GO+jjWV01RY5
Tasxq3llTTFKtpO5WhXXkUfwUEo9ybVlm3YmqB0XPWoi3vv5BtsHfVCiKbMx8Nau2i0roEBSYkUD
H0Zk0uP3qYCQ3o7AR8EDIHm6xFB3fwCL/dcDpPoDoDMFuaZBrTGmTygxQfAChszO9J+Mvuz9S/Ig
IwyioTPC5pLH9bdVP/55af351INRCdZYNYNUibfG5arVxuBTObi4PrCXF+CEvQBEJeUUBF22nYs4
1DQfcfTSuRAcDZWKkvnv7nVi6F/V6KXzO/R9pcdW2wzr1t4Z59Y59aSlx7JGO57wivuYL52H3VJo
p8uyo6xeKH2us/6Nbdm0aYJBgl11LrldMoUf8BMKdcnlMeO2SVcTdM0wh0TH5cpYPRxxxlAc91FY
GYj6iqRh4g+2DjM+/KddBM2sn36DFhi/YCUcMEJO+PFFkkVmB8EZNGaHGzodLGoZxyXwXrEHNhWF
XXChE3ypMpP0rlm751Hp5/DrvDZpBge1PHOwZ97+gZjPQR7626GWwBkZLsXxzkKh4PGeLKWTFOuG
LsHHYaiJz/Ma343tvTnKELDt6PvXIehiRkwHGXRN7rT2LDkpvuF5CGwWZRK0KRGbuU0x5JTcL7yq
cdeiU/bmkEKEkkOd4piIPoE6EEltBDViZLH3bqpSyvorS6A5ntDKJK8BjZ2voJW2jUeibPFXJjBx
nF88PHzthaS3FGWnKfCk7Vwb5sxYWRk/O3XynvXD3A6ua7ay/O/we1+oado5yZxmSSREXOASU43K
eiwrBqMkgeJJ2QVMxl3FDZThy4XsJ38P4arQs57K2XIzlQgz5z+SwGFybhuc1tVzPaSdtYtH45ts
t+FkkvKXKHIX+hLzD8QQunh9ZmKrUJH6QywI/cTOHYP0iFzxFhwmmWwgBn9x3lcfLzO1Wn/3WzOd
1OkUMrosAiKPfVPMJy3ySFDHvr21nJjcK8CRwK75DgYuq7Pa5X83MHYbCPmerii3aeanoDCbLT7j
hfQ40Cn55QZ66tNLUiRMXHrcxbqvc1ZFfyFcBsiWrPqNayhVuzkPnAYpnYOwHgdJA7oug0hQ2gzF
G2GzGuxFcRp4N7tKNFBPveaqfKceAJ0sryUep0VuRyt7slHBXbjSs9TJxi3A7+BeRG7ALviaBdfn
wpNPTwlJBjxkobS1JMdIxUsn9tSmGBvvBGb+SS9LstA04KoJG7k0wTuTbSW/Qcy7bNgeODxIacWZ
0VE2emC4DAp88qJohQUpY9NXU4HWUHvHKf8JWJ4gD8/5t3G+ojIS1UcEHZL2FpQoWBKfaCMgNFB2
trJvYRZ9HB3SRLAhVqVjykYyuB2rN73tljcPK8Qvs3iAvo2G7m/pKj3nJOY4xadWS1QNnrVCsiQt
sTMU2vayMXiVmwB+n4FuVAa1cRI6S/55AyjOeuRJkWm2QqQkoV9BAaAjXUmdAb1rnkSaz0Q+nk5R
Uyz5gWdFnDNIowf9pmXR+ZSm7L+E7ri/C3P5MZzyGRAj5GsECAWCEAxmsT8W8EDferQXdqViuKVv
N7LJXBpu4/z9omAiJRtT725P7xuuN/EYemy3K20gZ/C2hs9Xf+WkjxmGKhgtWjX6hXWKoHZQNm++
3GeFUVzwBf3PoyCKDqIYkkKscnqAkp6kVAGZUSb+OZ5QCTckPuoR21Vu854IDE3R/0nYbZ5km2t3
zIVkWB4v8VwCpospggborJQXbuhsmVQvlTqrERe6T78wLdFAYHdravf2NNzXZhn8lQG3nYsEBAoS
BQWan01WyZDljxxoRn4eHhIMBMeZSMeS+osQDpyau9AQI/LtMdh12fFBhMd070GbcBb0SDQ2C02C
JIcWjOQ+0CNQh+YVc1qi1qsP8suo3Z38YyX6tB24ofByUAgjdqyrCGK57jVwL5NslHUUbE+vkw+J
7IrSCijx5YhYYu/1pjLiEy/WNjCvJ1GYSKwG6NUbxmhVxjS6c30tNjE77kcHsDha6JwTTfH2I91T
nqyKYm8kAUvntQBQ0RXeeIFxrNcGVbMAksyWnLyvWDKgHkksGDEAxFnwcN5BfKOlkgYob2AUHfqP
1w4+Fjb9ujMHtcpr5rBO8VR1F3pjM5va47cVjhgJwVc/L1rJcCtF6nHzb/zyhH23lvvrqtTZMwPX
f+s0SKAjAS2J8/gCqAy5fW1i08wyYCxdHsysTaO6OxHNKoNJG9JbdZd4Km4n2rha6ZgPfjmeTJC9
zqhgb/GcPLhgkjfk2x8F48qyu05SYodSFLi3UwVkMp4iYIQm5d5Cg8t9Q1gTY1JP7/r8dQsfbFIk
k7+mNNh6N+OF0X7YsJzusezM8PMXkBJt2n+SD48NBvIo/qQ6Fgfej8QwaayJckllNE2lLNS5e7PG
LVyPe+AHHelPIijzyZ3iAiUdCJpQ6RrzO4ZsCV4N1uLy5vOgU0yLs4UDEofqpfxKNY/N/9zMVd5W
wJ36QTr59nI3p2P2SsfYMBI+eI8PFb7EGqkQai6kJFLyDy66/sxXu2mTEvBUrDUo8oYgj0Ay1Qrz
doI5a98tpuflFFTKIhnCwFCWIK8Sp9Mb9vH8Ja+IN3ohjG7PF3QRGC4FRwsiPvvUOn4ZliKu1u1U
qJHM7s/oIJKQtrfNRiKgwIZWu27t+XEoLmbM6AzS7VcajivYIIEdVndhBQuYl6mmxM9rqOKEtAuV
BNuL9Cb4lBkieiyaN6F2cAjmbBMO/F7Cbo23UyZwaW0R2H0CyVl06ca3p2uPSb2YuhiEIXgYkDlN
/HnevykCo4Ee0/r4YJnDabvIuP7wT+DJjGNxPYRc48rl4iydUOp80k/gJzdV8MR0uEXHJkEwxYPJ
sGwrMhuH3A8tGTVoG8G9MZffGP/j1PZCF83WgYdZHjSTA270n/kRhPetphrfn6Q1Hfqzln9Wpdgv
HryZZqOtyA0roUl5l9Y2fvYQ9ROQSi5211sZaSuYe4qcGsYEeMw6BqJHPWMPoXKBWaFQVve7p0O2
XNMgrIRUsNep/Xu0IT4Kwi8Vv3YCMzVWP7uxdjDPH7zSi6sfMaXDtHOGOdcsY7wfMLKkdU/NhKTV
43rqNCFPS3FFXrLhd2XOwKzz2D/JvjUTytGO8hT2vAUQYm7Li8MgRfeg1RZ+m3LaGLCZq5Vcy2qQ
8l+QHReYtIvklxOj+C4W1kIetWthPRx768zh48qySxV2oAHSYYXUUTGexUCsRKA/ihn3dlrIDagd
nNqiZaU2YQVl7QfgdRJbwffxIPL4aEO4iU2ETh3VL0Uk4uXDh5qshtCVWFztCmoR6xiQgKGm4Zhx
+NNLkQ5Z5f1t1XogC4yxH5aDbFrgFSZLowfdb1oYIvnNhWgMfx757cytIh3MaBUNSLy0Q2qhMNHv
bheFAe3F7fZMsGvZL+jh2K2HBmWG/chdt9ctzDzPmIA0Wckdo9ZUtziuFUzYye33zzyyMt596q0t
Wc+iuO06U4jbu4qPZmswogTM/CyXMknJQXI2wZfBoBV0SiZpD4rIHgW0/wT6FuaiV+/V2FoYDVa8
4jljPB8E18/i13DGhr9SS6rwIOAU0Qof0GI9VugrOmFg0uc+Vpiym1y5wTRM2Y3zCJLjIAZGfT0Z
q0MzPJiJXsYlIhy3WjrzKPjkRd1sBHawB8SNY5J+TtGyz/eD6/Qn5V+MFsuYVrC4Xq/hnXKN1a3a
4Va9DTSI6gwl5a/iiCP27b8bG7Z/rWWszZKyrdwvQX1F33t9lCjA6A6+jQkylO1vTdSNJidP1Saw
o4dNeD9A88usZ7kLmDoXdVYqm9iOSgjOp+E9k9W5OZfvKCEPW8TBGZqDSl3opOd7+0MM4HOFCo/j
OTO/55M6Br6pOFBYvKQw4aOhmf1PEtfMGzKgemhHlDb/ksuS/nRnOzc+rmvJtFw9HrAszkUJJr4p
ByEaTNHLiEwDsAFMID6X3vMtHvvCMwPqP+nsG0fry7D+s7zscKAL/YK3F+7zZlXl3pIV6AVwOUBw
MgMEzS6egfyZ7CE72L/OsT4qZs0GExcNOQcey8reJ4WcFGwdrROXUErqlgu12qP6oRp695NnNOty
G4DoRRPTdkZ8ikdemPPaUBgEpkXrqCeHKrU8L7vLVd3LwQaJroPIKh2vQLSlcSnhah6WIK0N+Vlv
xrQkYJWchS6wSmK9odxAwg8wSF6/U0FRigKzv8b50wzVgAQz7AphO2OzZQ1PoK7tTYAZyn6uWuCh
rwxV05uwbEl7PGo3dKa/VRkncZeKnDlBNtcSu9ygdGsZ12OXWjnoge7Z3Olq/fC4yprgkOYXxr1V
OoqyavdSVBIqR+cYXpvnG+U48sDXyhXF5/331tOEgIeVPf9Dsrgt7Q25yyNfUxHUFBxqqVwj5hYe
zPc0sunFpwYGQNV0zAhbOQu/keeyNOpQW91YtH7c/HeKU/W0um5agvPNeb8bxyCRA74cDr3Syb/e
vB7DDOo02gLDpus1Jhe62tTFg9SV10GO0zR6Y2eCkP3cGf7af58w1/WLprDdO8v3oRICQ2ySBejR
gSfCvmRh1bvgL68JqD9hkjVO4iBE7c/0Yy6HYfvK6Xex50+bQ2UN+8mhWGKdusmViONfuefXSiq4
JbZuHQ6FJ+cSOS72hrZNiU2EkGIOdeWzFFBY5w4qUpkuwTHG+l2JnaG2tnw5b6o2+1k6D4KAjWbi
xRRaM/GIByQfk4OOtZxaD0ul4kAIpoOlbdFRxARPCIJR2xIIbnQvhsB5yWhxpKlaT0IRj1VNiT99
3+l9/296P5M6aO0wsYoMoza/5315HaswfVVyqeAuyLGF1eBXlN93CUV9pYB7er1vxC93R+EbJo0w
Zx6Lv1DTAsBvHuzZYe3gdTiyWE/TiqBjMcydDTq9sPYZRF4Gr0Kn68ZpTZoQmPv19jzvVP/WRvDl
/sesu/rKWYU0ZbCXX1qxAbIc3IEh1KC58iXlZnttHQ10Re8DgiTuEX9ThgalXjN/ph2S9CTfH74x
C2FFxoxXTrZYJhNjVee6B3WetBc+Ny4YGPaOpN3O0yZ5VULw+IJvoCyV3UnIJvcX/W1D75zJfL5V
dKbP3LYHF2A6sYAfWL8vuDTtT8gLFOYgkIMWH90mQNVbRvoJO3cY5HR9zjN9yu495p8z6O3Ke2O2
xYn6VcXMblfd4zMSby+Rzl1OZX36kfR7wpl6vckl9XBwpDxCwBjE915p2FHjKzhTQeaxnniXx+VW
z5hJg3oHhBujSC/bmEesNsYxSjOlZ+8NKWzpQmf4bCGkwS9+SSccfx+g0Vjv4LGfCUKCyfq1DnB6
X3A19qm2/kpbSlxiyyz7F+OwPjUlYeG4t9pn8AauSeUwLqRb1YPf435DOaSPT+H5gdedjXYeGJTK
+PWGW8zAhT6r/i0d293GICaLY10hPGXfZvOm237/TM+xb2qDz0NknuZ/Rz5qL7AyxgblbBPDyfvV
fQxxo0a17v441+4dRAJQQf0jU9G7iSi+g46Ddl4gJtpgKVlexpMVvcErsCdnDjbGMuX0HsVdd/tH
cIbB+/27WuIpI5HWDV6rbq+ArG0L9KYvOiYFLPCxo/BiIGrKfaXMYlkayKzSdx9iUfXD+EiSj5Yd
KDTLLLAV4GOwuj1KRklP3dxqLBRC8xoG4zXgp5JXbG4Qo4YPNWhWbzjz8pn/8KFJF7WTsH4f/lGJ
mYfIo3V3/w6Amq/ZnGhx8H67ob6sFy0+7Jb7lUAsCiDrK5KnuhIzfv6iPqI/ycc4DZp812Xbch7z
dkCcpyZbqDdlvXospSJdPYPw0H1y4sAfq/ypA29cka4GEKEsXcxum9e8EbIobIlGYQGogkrXoU7n
KOzTXpJFEngbLNxAPnmDydKmYSGR7qZKFnf01cguDR94ZRmHAHslXLNLBxgd+1UfhYU9FZt7uf9Q
Vh2hFHVve/ImfLzOUMZI3zYD0INXB0J94VUC06JDh4By0LYja0iHf83yxOh6QJHCJSrpjjsLdC4P
kvtYumkFnymmhr5De7ZHnaczaL876kb+LeWbxt4yOSa7tESRplhnqFQI8gssG5rj6zf5jAcVCPa4
MOSlVMNIy6hVZ8TOx5o2qVGA3cBVM+M7XdMW2RgZcnHa0MBa+m79jwGGcTNOvjUq7K+g2e15ZyuC
Lq/x0fuRWeHAlpe++ImGFCjJF4UgeYxQRVPyBi2MhcoBP9fT+P/7kjjuJeEsfKtUBO47rDKPowHw
C43fsb6IQ5eoGkgDFjCCCJLEII8UlWTPTA+IxZNN4awZvJ5m8+EEZi6bzln0YOLMPrQiqFX72RDv
s3tLY/XrZkOWZNzGtmHR9Hb6G2BglGyeF43tPaGki3A6EasZNp8zoUU83TSbbI7FbdrMM3wdfU7G
76VjfbalTQRuiUNTSOvtXpxZIFoS/cpJPcfspFAbJVIrpjIjDrrLgPicGa85UftVAW4nw6m/CsrN
80FgaT1+ZZRTz+Nmzq326eNvK/Z1p4zDVT3poUJaRExxRLR6pnTc/YklpQg0ahS4T2jJe3c4HfXF
nYNPY1yWe/yBLGASnkXwMmdFLjUTfzjGnYGTmctHESLRYcZtQUCzMLng9lz97TCFuH3b7X037rTU
cPH6XbuK+zfvz0FDjStxD0J1OHZVtMzyspKl/wfJaBDUJP4JCTENAJbo856FERQe+dEddWydzyWk
8eF5Lb095JdJzDuKoZuYs7PEzX1zUuHg0pqkDqbB7TmkfLXPLQvFr4VksJj4YYh7rIr3X7XJYCwb
hNKFah35LFoFQYCd9Jt+eJk9FNP97Ln3tc8Mn/Y5lMQC3LwIjiMlTvJlTcs2jyTdPThGibo95wlV
RahCs7cUunYFfD7mjebY8ikHxrEqmD9S6G9c5ePGODwBdnIxZpxilHcDTdng8NpwynXjtsoSi8/v
ovCO9ns1/mId7TRi51VuCSL0DEatQOe0BGz0t6Ck7pQzz8UDwWJksvurXh1+EMmMTMxpXMD3MLyQ
SdBs1snooAJlSF96zPMofNN2es7uZ6XhEFBCYC2N4GuBjCLFHdJHepfA3MjrgkxXwkW8bB773GDa
LIMNJ6lBHLSrsWCqR4uaP8Q9bzBA9dNQH3P2b+JWV5pL7b4qKWer0xiu1sBlT8QQmCf1TuqEUbwV
JsuaeAgs74juWgSz9VfU9laopNh18PsMIgHdPseFNTz2WesnjmVnio3MrriBpuIaDrKKU2z6o9NQ
HRTWVjWNTKD5rS9kGy4UvPpfpZ94vVRAfvRltEfhGWkLiUprVHgVUSUFI7Q4TEIbr2pMM8P3dGYa
3EeouJaPy6Qcl6VY1jV7NJ6NpU5/Qu9Ebg9MRu2SsJNyUkak4dss7FwvK2p2hySIYkOLCTFZ9Ze/
WUl+1d5x7goB9CXRWYr3QmZsdFbk8rtnjHecZSs84CeJQ5E0gKf3+6JFg20XwdAscDJ7gd8uDa4t
aiT5R70Gto4mcgVb9eFBcZowLNJMEaiyfx8XhlQx0LNiTPYOuxDSp9ncc2W88W6iRMxIprvZeS5n
f+GiuoQw1Do//syzJFlWDWKyXOMWuEDrCqKoCtnEC+Zs91/fI0Q2YziR0IrKo+i6PzqWjpwuDv5a
N2R2Rhjs4dBxh8wT8Z4O/YnQx2bGkKEUu6gT0uzkpIYx0YzJO5RwE5HN+pKjRueIuP0wUjwGOnUG
qOSu0xYKYxFk6WMl+cBOd0KaDbgwI+MTv93wgOhbkmD3BNQ+N2Y5ypTfk0OH3yef+Svm6oD43ChG
V5BP0ZAhDio4mFrtT/4tnQQIkpUuf6FF1T+Fty2T4X8vyJ2F32jdpuL0Sc+PmMUczFR3PPSqkxOS
Pw2kNolCx5kAIsKWptzsjcoxbP/D/aA1M9AoPQa6QmWrwy6GF483qDgy9bztFnmCOMxpmzNSHJpt
2o4rmmOKJ1Y2IaoSrMwK+n2pfDiBuQVoLbSAHk0lvqkEi7+i05VvLF236GgfoauVZQJkhxzfQz6e
TkRY2lAmyCZLF2t5QW1fvOv26yTOP1pQM4dAdGD4g1wRpCoLmVj4lxnZu6pllZrTXtyv73gnjfxj
dCNwTSWOmyGXUVhfU5A3dyEJtNzTG8ccc1RAPUnQYbaowMsM4sm/FLjMd5zsfLcQAIJ4H/j8yubk
ayjnqA7L75e8prZ71s3xviLu31TnhXcaY99n4ETywfnSBX3JboazN98uiwJTx6A0TlqBXchDrJhi
YqiEGOId8wzsCi6ANFg8eQFMUCXI9+p9E1BuLXMCSOjZRFq+/82K9lRxJV0JXEMKytM/kr2KUIKt
MYeJoTHsv5Vr+7iobMQ/lelSP0IIG9U4meFRGYDFDsT/ek6+V/uj8J2uTTXf4wdXk6UsENzJu8K6
69pq5rmXikU2FELELd42GYjsTPJI752oXMQYbdaQnwWrvom0Y4FqUhNZGG9oqUDixXDgL6+oAqco
X/dDTrYciVsxcY5xIZgod41Mj80BXQhXV6/AUs8Pot5seAnCXm+Oflk/NhqyMVzoqpsjcOZsUJ96
sTyDGUZj7q6Ct2LceImFMpyItx+2bFKKwRzvV6TAbVim9R6PgBJG1WIxEvIesDyrjEtX5MFPUZ0r
QNZgHM0CRUCHSZ5Gt5co4mKY7sQSY4qDB5kqMyZ3ba3D9EiqT+HSaHSnwBXcwCDeLZC8t3NRYCCw
PIfb+0r7/+LM5u8AM/4OKIfmbvB+x1a3Efcls/72Reghbc26RZsHLGdFucaGA/UccuaOno6uSVnv
WRzL+07bvKuv/QKHp2CSQxHx1LAu2O/qeFeYD1KU0D0773BQccvk+kV3Dy2dpM2x8VoU84hMeANB
WoYQo3bB4rZv295fVIimX9TNcP5+nQrrCJyC/vuThH5drILUWPyyjDwcP8+AcFlPegXhQE9hXCXx
BfeUOdzalnT1183gdkvntF0kY6JK06TsfUODb9GA/YZ9ItB1ni8BudCQs08nQxrMztzxawmX5gP1
CdpB6QwhyWRs878JT+cgolbthlHiShopb1gROClX6uQNpzVo8c2UWIzyCvryR7fU6eyo1QgD+vpz
D4QIUUPRQh8Uez43kVtE2meOceZIg4DrWQu9o6ZJz0aePP9AMPaUEQM7KmHqJsj7tgWKwlPBiKUj
DmVMq4PEn3IJ6lAhqthBBTY/N0HiWfW8dJobBWFZ3/h0jrE1TaCh+gOqPmQGzS/dXMQSjSl98BVQ
ZtVbZpCkf3ZNxBxCkPnt9eAQjVq/ZuL7zupRlVamp8z5+i9KQjQOF3DLyYybY3497r8Cg+BsVL3G
MR5cczrFl6aaY382sH7zorr0IkR/NsYc9OsbDPXfXuGpSC7IqZ/woLIDTEk9JT7wtlJ4AMousvi0
WA9UBd0QKrmNWfFI54IERTLJ6CCEM47C0P2g9PQXYeiWkEnQkQacwcAhadQanJPts056t0oT8IEU
FYanY+Drp+3wGF72V5hCmOYGqxgmhHPzo83UzOIFq658rwHbBkA5JVDPoyBmSnrDARGYf6n19DJ5
b3dVd7CtSs82j5BcIOyhfhbU4lxsb6fs/IXMr/hNrtP1KMHsBUH6DOXYNrIiUIBshoTAERb8bTio
QDlAiP2qyTamIDXVpjUw8VHctTJY4UoF3lYYvdY6zXjQ2wcpI5dleJfqTT+J4GAgSwfuAqQHK8Oj
N3x8DnPAFGDNGSGsOtHIqs/Bi0fJOAA6OyG5qlUC/O2wANiN71Ip0o0ohHwl+CDTzpmi+Q7k2h8E
HERlDUNn63ai58PVTazbn7QrMGQAISzoAeco2a9S90q0FpDQ7xQKwSzphwlCu2egbAdRlP02xs++
YrvPePwiInFVtrhVpI+H2Ii4Vv8GmoSN1ClIxGEEP6Q4DZFhKBkblpWR4rGU7LpxzCt1ECV9Ppsp
PfLmnof2JYMR8P1DGIPnXZ13Ey6YhAflC3t//tqhqpfDFl1iK0WiQfYbGWiumYN3KnDwe69+mprV
wVCVXhN7k6vm4EpnrQFrb6WBVATtsjKnH5SXxG8AkZ/2ngQsjjzeK5mivJ2kAAqneIKT22VfXQGa
c58ZTYkNUpiGux6VVdFMOpKzj/Rcb2QB++MLm0V0uMyJcuLmuJ+cnFbvipdXaGneAK/vmnHDlwYg
36FfpIfsWr/n86CCsne5MiU41GtrfI8HGSzJDaTSCb7xtrfjbKDsuKK6t0eKwjVqkmQXSFMyWtEk
EHurzqLpIpenuK6E52/6IRBed7tQ9ZZLCs2wWv8xUYes9ktniVrqW2MJLwMx6bfHek+QQqKEHQ/E
F7lBgltLTOExf6nV68YBoFU+oAbRmx/4v6+50GhMJFRa+nYOVqd5tiqq4LhyBbEu6ubWtlaCjMTz
NRiuaEy8sgX4G+Mrma1tZlFlB3+OR8lAr7LdFSmCYaGQBrfIzpMbvTRNnG9aI1uoxQJ+cdRpq0mU
v4ppUnfFG70LU4Y2efHWeJOYL8ucHUoA0sT5LA8VJVHg9EaGTCD/IeW3vsrzn+7IGNGtKnQ8qlx+
3qk++DtVev9ud8YWp9HmArEEhRa+lA4rAHeFAW5MadHbS9X9p2Y51w8NWx4sWFmmYzcPgzzS4jKa
Qza1mEEeS5YgE56N7DPoQrE7Vk7naOfB0omyVMKg4i/vORN6970qefWyhVhC4V0gs2naUGAXzSgE
lFQx13TeLgqfw5aXzgeZS0bE1gMMS9ozXSltVx+/0PeTnuvSfRAKe5zGp2iYuEJE/s4KK92tKBp8
FG6nAswIde+4XhmhNlRgRnuc9Fnl1AboymZSLgCpikhJq3D0QRNIsbYItpfMsln6IAgDo7zx9osW
LdCE+ejhWFjJ8LgH6CNKNIGmI2VOpjQTMhDAwdRu+3G14ZfVQaMKNodUkBtsvFZLuxmhY9ORr+5t
G/pC2GMMZXqtQSConleGT+sMi5bCFBoaCgcHgzQmxdix4nHphUMVDY0f/D6F87E1867Yt1Lq35t2
Cq7aOjKOsPwuXC3VP9U2MJ6S7c+22cXcEehK/irEuZLntwdHyHF2KjS56cDdEp6wZlYEK2I5fEM4
t3/YmgFu96FMRn/f7foNk55Obs6GSxHUc45lvUNnR8Df/ierSGvnY5Nlkc81ja+UmZGZcguF6iEa
wSMj7672aqptKxgmMWIft5mFuzBVMP8Xez9s8RYvvo/Zn6T90ZCLMLL48hLAmWgBbPGeWJ1eBQo2
n7WdG1FtVTrIKcjaLra5OBr+JIS3c9uej6m8YO8jPNprpnpSghVrlmJ/X0kdat3DDSlZUfgfobKJ
EH68R0aHwqPZTMfzqzuHXqwzEUcRGOBMMfMja9cKFNFX3DwJyyiIsZmOGqidAYlr7TticK8DedeW
bwdNu6n90qaWVmsvc02vy9tGVZEvYnttWaUKIfJACwLd+hF1v3knu5EoueC+0Kx/2bNE96SVmZRd
ykvHKrSZM4sjy4KnuLGz5Tw7eJZmku8u8ps2NPvbXU2oDp57OCC+U37JrvultONYEiZDd/518KH4
Wm8xHgjvMFHOYZSkyYU9jTgS1L5xtwJle8pXVD7iygwzwKiIIOwmzMxQYljm7brcMTZf6GSM5la2
Z4iUsHYR/OS8UZouBKdXK2JOjwdMsrAGAbGbuC0H/wnpQ/12ZxMaWUtLRL5g0Yr13O5C03ClOnHZ
Mj2sdw/W5rokfFyd3gWTm31zHJ66CaLktWONES1vzE1izct/mVBvwjkceyTk/knzD7H9rI9qsuaF
V0Eqp+EfU7ZGyfgdUJDJ7Tj9Ga31CuFlvqFPmJEFc0gz7l+Kitlee/BXeSlHU/UL5NErgz2rxKwa
6rnsJTgt6EvzSTQzIg0VjDUURfOd4+3yjaxdye5ymDE08kPmRIoj7j4dTdG1B07pFFRXS/fYW1ik
r4ONwAexIktX/hgs/8gHDb/m+P5hldObDJrm60PR5Sw70U3u9+6cznZHmGwPMxFFpUfsVkorKd4L
LqJSRm7kgg+8W7ohdp6RMTEjoBJBTxO8UqIzV9pk3dDo3vOgiao8eE+UVWpfbqdQpPZi3a6p7Y3S
nbnJyuequVfedq5abU6eev4X7mC0bsaIu7XR3l9eZ+0BoL0TrS34tUwcrcVZX6nPO3BegGWhrpOi
TZ/46A792caEydE6hc84EirzKva8wSv/WqGaMzYIW8pCDt0ZgzmCngRpROJ6VC+gU2uwHLyQtemD
dLw3m0L/2o/Z7V7oodtojWgKFV8t3bnxYXDVwiaquD2OjVoq3aLd+TiQE+Rlo2x1PcmC0oTVn/4z
BWWsfNc384nsmN8gUmC6c4HRH05Qd7ATivmbfjD3AWZZeOO86EozivdHHH7I6+VdWaLxAbxaO2rj
jUtZPf7NP0X5Si6ViON+7DoNHwy3wmRCZoGc37habvmrskllU+4ilFJYN+xc8XnLXkGG6AXTRvte
hF+jNtmfc2y4l9lgvGwtX8UhwQtD7DEnKcSWZFaP64j+x2Jt0qktxV9fGXlKmcuti4DxFoQzWDbc
b9L2C8qW1B26c88sIFmt3ttn0jNqgZovd7egoXsxJnP6DdfIdA+yWy+zkTqfufHZ5f/S/iAmRarH
0PAOdR/eI1bTQe/V9D6B+DpmNgbr5sPYOJvfEkbjKIcVxGHVj1YBCnaydqBMaAVJzTAbbELabt6f
2wtp+NqbzCiBY/Xn6GIO7NnOtoTg1ZE8IeEdCLXsT327nF3xZn+QBOxXwzFGPFlJJ8NtroGz9Eqv
v+2v1Ci73qZiuxAU226zvNg6s4txTxUCKg6VMf0F2PZ1G6NpOxjOaQpOe/Ur20o8IWva5/it54ss
8/H8076xhrb/S6jTsvjSgL4TDrSnRAW1dWg7FYXPO5/mzgI8f3Opw6zTw8pfE6BO6G0JoyqJoeVi
IWsdmlTtVceSM3CxyKf3+m3BLIPhQLi+DigCYvR3rLq58pEHJ7FfIY5bel2oLIxqr4GFVciJosmI
pnlyvuqEjfwG9ntergBO3QhNvcX8PS6wHqWDlVolYtPNgnYv3M+LUlbbVanVgK1Dmi+EIkNXPeKJ
GHZC9KRdlN/V6Hs9Q49RwcdJvMZwtCaf1wUL4UPSkmgws3L21vJp1cj5rTaxX6eptg5ELvWltwMe
/Q/PNwUXNiPVWaV64/RWbNmOK3elP67yFlF8s0bZukkAfddMH+fIw8BnpdiWo0k2N/0Bd8VnJ4iC
Bp1mdpgmNSvtq+KCi7UiRJyhA2q+cEKQSGwH1R46Z6Q+Pzp6meLOXC5dXu4iQGyEA54UikcESiCE
inQt5dXQA4YwCz7VLRwl2+I7iE0UkGN1bYW+TrFSHsKFmbdNsE6KM+1UEG3K0MT/jvYgXWB1ZSnR
IsYqbCHSWb5ILN23euBEAc9cULq/tVhd+35Sc5XUzC8qkIHaIhjlR0zL0sOKIHvNCvfT7vB8k62v
Rjvcdc52PeC2BDmDCx+BMf9rrixZtKT8Hu76yGFa624v9JohOGh1OOv2de6auRpyh8fWFlCg+by1
TIjYOxl2S7yAUtieLP3102AnigYIQgEG+igYYGdbLayQsvkpifDbOzE9n6drUtzwfmkfevaxbSqt
FtOvcfeTjKoNTZNbBOe4rViZczU/aWpkirMn7uql3ycVPZQHXKbZ1KCrSyzh95nnXGPVcHHKlfvx
w0NIZP03WNVWGD1oyBl7PV5npMZHqXiXnIqBLT7giytAL+B+VjXjJqbt5DOcqsgGXMfTWUgFeui0
hWOoqsGHiCPSiiPEFr14DtM4fAzxs4kXiIu6/Se6Nf1WvTWzZ97s9A4ppFl38KVSmfK5tOKAmFB/
+JMSH4DuCOGcEzXGtBmuNxEO9wphOfLNq7yuAEHmfdMiMokxucI/Wxmgb3hwCJmos0ki2nvPhBcq
4XXLML1980FeRLndO9ulFyHWXh0KuhNK1ZX2a80H19ofk2FYJNuuwc2Q9IvpFYJj0SrodHNhBKrY
/x3nK+mKJ7nTXpRV41xmP+4x06Fasc+DSMSOglSudBJjd8DYgMhy453wcsaYDURlxH0LKUA7MgDM
wm9ah5sarXCuf0sZZs9LPWKUgJ1+6oQyPNlOEvhSeXrxlUOZF8yMMooyQpULNuhpsXYbYC2KN5sJ
3QjIRzfVHSFC5phDOoDJ0eHTElIKuLSA1u5NSaT3+yASUWPjHj8UxIO+wRJ7u2UtoIjXfNrQxwQ6
CDq0yc3zRN6n9sbOR3e+swE3EnjAGF6LCRPRIhL/3MbtB6OaeCRoUc4rWqFHGn+fpKjBcFrmj4ek
Dv2EnvMoCjhHfKFk+lwad1ft9oJ7Jk6/pQsZuD582kuqTd9eaxf62GOtvCVD2SiwqXGhPxoFMa0r
I5VAZ/EcVmus1o7I/spOXDLFJLtA35hklK/dZOVrgSxrD60EVcS7MNOOg28SQbkEagiZ9HOrSnXV
MJVqxzkYDzoF268KIpgeXhvNvIjMg6oVu3ikwIFC+B+2Qn40XCQXLWpgGMn94KfdgtCpvYGSChvg
fafhBTxvgpRzj7T1XKkZ3B4Kg8F6Mz4orz2gY+jmihdbjN4CFLYMAGonlOakbJ8H8uml+JceLAQa
3HZ4QqWHf/f6hu6QxbuN7SOpX8jVex8JqSEnUWY9f3WxWl7A+uPREPjxEvuiJCrA9YTJ2uxf35qw
3t0AFBUlkHmgigtxawKJ3I90+Dkk9Dni6WthDQ2Z0yaaciED3Kv5TG5/fxkgWsRNuY6OpL7ip1Q/
OQHh2MXn/XR/mmgvfae7I/7goxI6DvrM/eQR3iGNiWKs9KdkwVLGD69TgyGTrbzjfq4YHgQFfl2O
MhsKmzNyuOZbgbOYcoKL9ZnQBhgO5YCeka/jXNEYAujbNXLjzGpsGTifpnk7F1sAG9D1UWwiuzQu
HClX3nQbglz6yhPJT3myPx9uDhdBtYxawxrk6QBlaIDwkQRe6ZptExrHilauoHCfP5PIdBdBPniy
FbKSi300kKLOqGy2ggpSD3nafJOdC7n9Qg6VOxR/YFLs6Beb93X39TMaDdZ57kW1evcQzH5xL567
2jY2VEV8a+ArenRbi9EqjPhVnsq99HRQ7oyNhNqpF3tpIfUPLhYq5u4Sq2pfDFqXISPuZ9/vrmT5
Y+eqQAsNM//91enmr4yrAPqwssNsvdlQbqJUccaiwia2w5uIa9dft+HZ8qIwMpD4j2tawmjdrxXD
0cvc4mnuZfxRhsbojX61+RWOyMI1K7RkS70zulYXlDq4g1fzGnQz+F/v9F1fXCC/kuzLNpnATRQE
JkHUSd7Qz3NfqsiTfNigivu+sUaJZ17cPVH26QjSXUV6G/J+M+a7lO6sgsbYjVAOcCldaqpdGEpI
zo9ZbvhLUiKlY8K5lfZTqJ/Bw8dgYOCZ+aYjkMC7ZHtQvTsrfXPxh3miqVqfwe9T7qj58C7O7O9L
bFODW9dk3SjiTiYGFPWKUOFM/ROgKiKr9acfM8VAAsUjLasYKe5OeZM7eL+JAW3SJpRwn6CO+L2c
OMEvOaWZlMJN4Jzcz2hXaFQxAE5DBGL/gLF0rvw4R6gtcYEVtIFh6B1ET6uJI37FcFevv4KzLVyq
UdNiMwIngoXnYTfMv+3NUOglO826XFQT/YhcFQb2jQKiCS4fOwLudtVBlVTAHlpXE/tzYxmItZTZ
2I5Qk3I1ba/Z39+PUGlg6Wwmly/I+U/LIEpRhrZo7M6wiRKX4wdN8HnLWhZuk58HpgZHaWGxEaJD
eu+0FZILpjmvzQbtA69QmqRyGRjTzWhHngG+5eOLDHxnfhDpAamZi60/TaAwX5dHyJp1tG5PjYmN
KrVbfrukPcX0lXQtbSkHIrv+rL3bUCSWtDh7qC7I2+N0jORX5gw3vxLNAE3kS4BBZJDQZtt3FMeZ
+NVOafwXNZLWBxHAEeuZSBsCWvHyd6UDAYN6S5zKNPZ55X1Ogkj+Ay/k+PaZcOpOLOU4ICuQW6Sg
MraTWx7MNn1Swh6BG5N+XJsbnbwNVNgWmQ9aaGnEjzNijswjXWByMFwiDG5GSj7IePpXF+mwoqkg
P9hHSUx7FZ3XyipfWl6+icENJBK8YdZD9PGLYKfMNPYF/tO9/dIjItjJb52l36pcYix2VL1M8j5F
K1XELwoHHVC//3opjuIaDrsocQ/uY0qofc9Tm4vy/gNtpK2UlKoiMrgNYl+07fYZCSBrczDEfBv7
bAFh9M/fQWuE0vNghIUrKOThgsOvEJpsCxOnUzqyB20Id/vrja9L0N86yNlydjD2USU70wFtsmhi
IXCTPu9wBPINtBs0os+or9vBURGy3EqY6PwVdxO987pew+CYHFJfV2DX2L/RRBniEseCkS9+fPnR
jbcAVsusYAgX2t+LVpVjc1Ddl82EZFSRVvjFJMP557G+uhZ8+Zm4sggeztnDDC46m352FuElNq3F
IyrOwUGjO6gMHhE9ft/A1xOxw7Lp62CaHZTQTD4s22o4WHpWFNUA2Tp2RdlQmj/mMLoHEaun0REv
K5whKdcwC+xofGEKEfWadoakNN/3UVrAc5okVPlQG5AyLW/LI5el7TYptyIKQ9w+UcEGmwEIpGsE
2brzOBvGUAk8A6Bu6HYWZItrXdkHOYZvzdGhbbJkozwKLhY2SFJ5J63n0ZAwBAz48SSxHAHJTQke
FG10aNkcvytZ9GQhOnmCWR2Ws7zdFg8EWOUhRc+B5u/GUvlqojmWZlG+A57NfqG2rA6aWdkuNr2c
tVc2/Xoj028oIEZEF146ivXWmedp5XZ8ePWxzQh5DeEuxhEe9QN+zBcC11rSqCb2IrT5LfyeufNU
ZvID7GAln20yXSStGDRCiiI87EH4ueUE+9VDcryd5Wko9Pb+VO1dWEK5HOMEjJou567qJ2Ocqr3b
hpLBQNE/ZHcK1lsibqcL47/OPQIhBEtlF7DeXskDqPpIPcSGqbPL715LtfcIx3sYR9NyeLxCx6HO
5WyX8FnaojxEgfpTxrpjurMsL8k5v3Crez/dTp51vqYAoWXA9CBjQOjTafJDO7q40E5CDcXXlDwX
FFiWgMG55MCzcdD1x6iEmn509LaU9h/F1+V9pm8JChDkmb88GIG9Ql3kzRTtuXYkPxM1ul7evVuw
D0H/osQCvYYifx1nPQWIWFpJ1AZCHCAb/IH4fZ5lcIpHTSZMRd5a3HfscL0sDoA3bf7OI+WWFihg
Qiu5uoeV1jtsq1xPII1J8cKGx3/YKXgg2gkuEGOoo1YGLDck31XWV0qyE4YmyaG9V5s0jtmKpCCt
bBRY5QnmpI2UsfVHbJyZcthg4BkoFgRtQhTICA8UPTubFs1Z1j8wd81jbsvLURSY5f3+9PrGTvka
2vxLOgfJGX/lOzTtFI/chGbSfc9H1YAqfmzLgj7/oXQ70ZQK8vnnTTX04CLtG50ucuHkpJ3b6j0E
Gdz1ZZc60pI5qQpPxf0TFF/L15FWW52A2zVhbyjwzyFd71IXdmm2zQGfh6aaprILPW0V7lEGbSGs
PyydUf6czhRDxolFq4c99fai2yEMCuVGJHk3byOFVG+twOgaHQksHk2yNkcw9ENa4wVqIZAQ5GiE
dZijrgcvtoafbkiSntyg7AgdjGgwU01ZYf9ZJYs4cM5Rng/A2++aFj50whxj9qcSUFh3T4d4YFkg
IV+iLBRUfzLNaR1xIccRX/9ldF6biZiW/05EtfjzLnPJ1xUKrdm3I8MDP5ZyIOgO8hFohD1BKS7D
O/qtjFPsQalgPDIZTgNTQ9/bJiaQrLDwBRQoKR42rF6Do9yiijw03gyYYsKJx3+Ul8o9lZk7Ui7u
Vstx6Jgi4NOZVwTHyyjhGB3vFvrGQhiUyZY6aqh/lWVFvy8CYYs0H2q7tCk8cgOlqYSj//sGDp4H
4+M2TdlNRALGVjTk1HzgYcyWHsEq7pqroiYRoWOkv2iFpivV+mS+GIY788PXn/YkjoLQTynsPtja
L6WZIoROCm/2kAmWMymFxOB9H8tPqrrM8kq4t1wVgcdJlf0S/GHu3ydvc7LjMKqA5CTBNe/7Hgdx
GENevVUAa9t/ibkVVo7XL8FDyeCRfTaUNE6ktmUcNF6eDkzS7l4vFJoqfPf2NuuxJJfH/+YTeCYl
5TQC+s3CMfe9BLIU4L2EZ872I1sYrSdNgFCMZTIemBle547QBT5ffLgsczPcnbnsE4PNNV57WCZa
V6hPPWsuP3DRFXPrFSVP561Tkr9nTREpGKew9VSPaU6xv1AXohjPC5LfixuHS4/weENI80jzCJbq
WAareoxhuEtdCscJI3A/AM9bUMpKdL6nTSvrkR8uqmc0ui3Z9UqNPwiVJkSdXXGpsEm9wqDYz7Cu
0FljFwFk2vvgW0eM2WiC/Tptxl+psECu0Net50WAs1BmuH3WYh9RA0gzUFVHpj/TXAmmvAVEgvYd
BqKZmda2BHjndzdLwXKtkeaIPb/1fDBSnzhdFXYTEjh8eg4HfhwKosWuwTqm/qiiLbwDU2YKMR9g
TmfZ5qhgpcLD/PeQ2r3/EnQCKFnwMggohA3QBj+CDa8IezOuJLLc2mAn2ieG9JLf8e250fauHGQK
j2iqnQK3tFrz1a1EIXcA3R7MbWhLZfNkY1ggJJvsM+ZHVEz4BHvIfAEFS6GlKq4RBFYhYgFeuMFG
aqXZZD0Hyl0zABgtX7mlSvzdTWcsGR0KhkoPNrzBlecrwXY4LbT62k8+oJmQpZDjkCMxlSEoxbLI
gSYA3KFHokzVZuCHCtGuqbL88wFJ7IpW3HAWyuM5AFALqP18b1ZCgD43RC9QDXqI1QMYpUEo4Nq3
gQssZCKPW+fU+I3rs/JehCWv7Ve0+5iUl0TCW3Qjh1Zk2MSZAUAQjDAfy42kfu2nv5ewIP18JOiz
KdXRkEF3RkqX/9uqRnk+aqcwzxrAJsqZqx94p5qI8m+4GQmoDak53+sF0F6pNlz4wGlxpdSHqP4h
tj7KJYzrsXiILSD0QUYiMiG+iQuLvyVVvs2BETVbX8QwVED+iF/i45FH1RCAzeNXZm15LDlq175e
aYRphmkGUM+NwOosjpli0QwkEOgqJxLJHlR+S9wIvV8eyi18GtB1iLAQslwQDUhTh/OU2NkEwLw4
jUMXv8rCLlPbSHZaG5w9GhYtbVPLKuBNgq3CesMxJqXDf3x/NnGv4cVjnxYF8NhU7mxbPhMhRoLr
TK1LnnCKzJur1U0h26+ADH7BeUVZ7nX3zzyd5nxKW2+jNFiNvWOplU+SePklMB8qAUXfMwxv3aN7
4QTziZeWXW9rI6ZflYbEaqhut+DCe9mYKVduD1fPaticW/djqmmyduEeIEvkqzDN0HhFmjKy74IE
Yp6/yn5LvP/lxLxHK9ocAcWSnWXknMoZKiYECydo4a3yUxnwWW0+GsWWGoQbwgITJJY2i5J0i4eo
7qUhYCwebaBu3l2xFoC68MDRnAWqgRC8+/6DT8DbVj5J/h0z71RYxo6HATE6RKN4fjMzOm02yWV/
MAz585Q3kCN84XkW8LcOkLBeJW+OUeO0E+0kHGPaQXEWto3YcU7nW6LwS12n+N5sQhAEOCpzwhcr
5XgkGRH+hBCvFzi4Mbor7hlOUXyKJwlGTtD3KOc169AWsjsXYKx92W5HuGSj1/PJB0qsepToQzaK
JOi+uGPIBi9imzNyqpaC277/DmsO0c80G0BE5LoVL7RAbgPYbEvoYMXcwCEWYN6uur51bpL9GNLE
ZnRbaqcekuqm8UnMsF08Dct2XTGQPetKCJ10WPSK+VMNzayV4EA5Txbe3jqR1rLW9jZjX7DGxF7P
0wxKx+nfAYXJ0M+UOgHilRI4MsKA/zhYxjbjNNig47VbMiSdY3ovtDyhyFrEKgEvGHcuqaprediE
Re8XJuXKQJ9GvezZto8lrQrR12SIiDuKDEvCdMatqPysE8g98/w/1Gg1ImZyOsVdtG5KzBTi5Q87
0PwELpSRiBIl8zXKqbm7NKXKEMMTdGyes+Wjj0e/G96I/jxjIw+RipHIq/tsIAHAZEzEwwFimJas
4Vx/HIZshX2ofNMhOIK/k5VCF8PiPAmjwQFtmgCVDRgXPi2wAFnGDuQN+vFzGQe1QTUGcOaPrf0E
k4IS3XUGKIQkxP13iFXF3uSYYVxgjBlmtVmhKodZXSXJXxk92SKoNl9UDQUwG7U2NuQonUTWXaPs
s8SMiQLB37zpUSQKIt3zGEZX4wu/19xxlpsvAuXTHXXo06vPAdrNK5HcWCy5DMy7gL3/11g1qcXv
wavysgS4tYgSd4fVNP/qjuOhQnFfyy21DFPY0vZQyGaNg5SiY/QXKUf7UmY2cJ8HrLdokpI1zN1w
ao8JZtaddO2wrqMXgyCyXzrBygk46a4pqPp3RKT3qNP8mNPf9Rzldc0QnBXqPDFWLiQ1e78l37Vl
DFAEY6JOI1kLO4WO6lLamvPk9ICaw1onQknXT8EJKyrEvBix7hJ4CUDAWyGURw7/i3TK/h5o3RVE
pUs39E4F9XQ9CxSwJcZuppUD3mVHAJxokH8cPNDzEvlhG+cRrbOIcysI6YJl/O7qumuSpuKAYqK2
NPf1vF+r4yHqG4fR6V67QdFSHHOuopxjyeBzW1hhWqZf/MG54g+VAXZid2UN5VoxG94GeOpvmNqo
ijBD13R1UG/WHffxRwEGKXsCQDtJsaMpwlsyRjuXBNSYn2F00rdwyeIdovse8ZMo0+E44A+A4cnF
GjkgmyDagTzcqJLYJ+z+RiB/ArLelgOoEq5Iqum9NydzwI2DMy/fE66ZW5rAQDn5n4xpF8nOphBK
aci8Y3DEk0YeO6fMu4QiffyTd57VNau4U2AUDzKQXdvJGKjICln5ENDR+Db/QjL1fGvjY8y0oypZ
YUe7BY1rNGxZYg/Bq1WVM79g/1VCyECs+1JgtFPw8jqsMHSqR3qXjDfKQAGflxsHBUywcvkyxpWd
32F0B8+oZByyTEHH1eRl6pX6SUkpAcmMKKwzaJ0xGMW98o4H64cxGbtsYbCqy6lg9ysNcEuVxLGl
Djh2RpKM5xn97oX8TKUtkBsOF3XG7jgfKq4tfKvmt0wBdMSqme0Y9Mo/zqHvYNr2KKET0nJZrODt
p/HNedXaRyEdhiiIlRl8C7Jrmn3DPof+QSEvp1Isbx+nOCVXk/9cS9cdrJ2/NxdRSl4Qwrq6vVHq
S9MKS+ywWHCO9Y3PElp4HSz9U61iazyPbBG9W3Cy+pjZV8nNOUsUUAcgihvPt8a0iMRCFWfTsHIP
u9kVKgRzMmV+d3pwISWOE/SsNgNg13lJ8aPoEjwiW6hIY7KR5jYZLzbFs7fw+m5TygETiOtkNQb0
G53hurvOTs7XfSME3LzJpcKOjJ3CvWaJOiVZ2oQLefc80ewbjSskHnqpGAdo187c52r62g7Cfa5A
e8Uf+ltgaEtNswYmQg5y9E3vrSV+xD6rPizO4fH/mRtPrz9II02rQ0odbiOWewa9pp9WQa9uBd5E
aFWlX7Xe9fy6IUgXNySZAifImz2ZuNv1LDtRRYGImznE4i0XumiJOA1TN54fJd1XH1IQ3aApGJnd
HKM9VdJnPyv94pVvlBm72Z/73MMjOWP8Nu7LJhG2qX+a74GwqrZkx540HXnk1XsSZL4msCbw4+ol
Kwm27HH2kyPMHp56qqj7LV1xoqwx225XrYN8kWRETvi5NP+agMS+WM5WaVKSps7Hby46V3O+faIx
aGfOGls43TGFgP0RACpkz27towUFH1dEhFVlf1Wjh/Hrsh/CByFGHhcWEXOWx7LIcOLtRzUpqlpb
0PosypvwwkHDbFCWVAIRjZB2Poj1VymMEy1JWJnahVej2wfm7hD8uiYN91ZVGh5FmaL6nNsUth9q
Sf6/E2hcHQ0g1ya5s1Z6onilpFPC+lEskYrVzA99zt6iXVWur6RVD6IcCiyxSorzIP4aSzc0UzcB
2Jp1uYiYkurP4NqDKgfKgcXbgpi64JJRbtOXaknSZDHz4gs5+Qdx1YUmfXr6lUlhBLiCtef6C4/X
pGNan7cp2zZGQaLbH4VfJ1YRhRy1cae2+RVAeENeSXklTL8NSZ/qMgG9uPgkE33GUOqaix35tdzk
NBO0Xjx7ttB5SoRsWX7iAI45MerPqF0nXGCQxXhfy2fheRcYWqZkAEd3LzVImNIJUuctP1AT36WW
Zfy1o2EUV6Nlw7jqMBlrIX772kL4c4b1aMVU5s57s8rtL4E+oMqQhwThaInoKPOvl+oMJbHlRBqf
MsfitkDm3aD54ljJKTpNrsnOE2jbvb9RdSv61o+UOcxZA5zj4iHPtdpIwL8GrCoE9oAcg4E8zyeM
TW3FXkt9I0WJjvwX9bgseRWjiUwRX14JeXnzjH+rIZgL/gkN6+WeSKRD4l9GQkFmKC8IzDdI6h7s
AFMJ1DvdJHgLkWeVmMY/XfbULxi03tXJRa4tTv877LqAiwSa9s3r/pnRafy8n9pixSFuzh3mdNng
SOQ5vJO/ebLpzKLvE98NBesuBF+39TIKthV+mPCY/+oCye5wxz1tGNjCxIAIg7I6m2QG4U/eZSjX
lAUHPn/+83UsVXTKPNRe5npN+Fbqz0XJfQIVC2PA3WTT7eFFIK3SpBcnjpz//iLkBwf3NoUqcZFy
s7NRBNzWoqA13gMjnjcMdY1NxAZADVe9s6FHeMaz55iolsCSi1A6iJh4ZUJyEuO9J3swv207+uj8
TRY1xPJOsNgZVNf6pUczpVAQaEs2Bin/sxdF5D+7iVFW6y6QYcKg6OSYDE6wIAATumhhXFAbRn6b
B+v+ssjt/dY9peuxyXeGkfty9Yu2nvaaUq/7YW5yEVT/5VIO9494xJXgpPw56uTmHrn5HLQwHglV
t41oxDZzMe/ACPHPBf7KbbDH/uTNys7so/ukZk8IvO6nQFLnqJyp9Ww2WyxhWb55dfK8gMlTmWIC
aFPkiDHf5RBa2b4/y6My9OJlr/qcxoMWmFePpSVNnIi4lgugMbCUtew4eqSlQdSS1jBj1JM78g0b
vGcunrBBalfkIyjRqmCupER5WO0BITcaQCnT2RKWK94EnxiTF4ersmrAqk+5PisIUoI/C1cs4w2/
EVFq4HrlbZALT1H+Y8wwiVqPU8ciE1Z1iNDCXEbi68ybWu5JpPhNzJom526BEwtIIQdF1i2ur001
t04t/Rp34jhn0cLQ05YXKKkH0p1ZPjsKfdJX41E332xCdkj4vVBU2z4dnEjFg2YgmJSf70RREFIW
rxklgroMW1Ud8feHueDHfsZaoyoWVhPc/r1SZ+XJ57sgDcoHFOXVZzfDpL0UGYwuU3kyD0PgeL3h
zcY8AbQvUBK/Eqy+VKCEoREMG0vUMQmDcnYj4V9ooR3sc31rF2Z/i34dweEySt3fNRZAPMWX3kwD
orCejAv90gKHpwP0oyD+eW97psmV8kwb46Jd/ox6EQFC6b6Bvks1URba1KgsM7tGs4YwMGLvNx+p
7CsJGQEh/OrMqqe5kjTlvzTBh0Y+39zmXihRprRUp94odfqQj6w0DeJsCgmp0NKESttT7JRmAW+N
7OkoNvUNMBxCLMZBy9NxVXhxiaYK/oJQgBuGh0hOZG9KbgUqqzP8bIFNEBU4g6jKddrUhmKkC5Cg
KzrEhxA3FfZcuGZI0hWi8s4s9x7JLeEN9EpuO9qby3FdtqUTGwiBhz18bqSQS/RCuUEJzXF1ONqY
2mWLhHAfr5o0pLKI6zsy0pLb7U5YcuoqzZnAmx+dYVa2++kleTlVDrBSjNmcWpGi3+KeBArkfFVC
Opx+IOZoWGINoodih+1Vu+RWpb1sSlHed1iaPg9FihbC4Xpu0TPLg2vgFORMRvbA93xyPt+x9EcQ
gAC+3lNvRzG5lYrMqW3VbyRLx5ulH7Cc3Na49imp7v2ZwlUBI4c1B1jAwPJSZceJD+0+NHI6S/m/
62M7848q8qynHDwVeC2kdeURs60rqcaAyMGbLYMG/EQ3CNFED/XxzPOac7876pIknJn5dykzQ4VN
7lwNVr8Fo2gfAh/rOfvFX+mmYZcEjTWI3yj60xhxgdjjKOekC/tPRYfhZbggeJLLa4sLbyxAuCbi
WthbOGnG/AonabQW/nPCM1U1w/z+HhoMa4KTN2WAIUG9eB1h0ZEWG06quKP0os8fZ9Vg15KRDrNK
2jGRwyy5w2d/1yQgdcRWgVW2M+ZZdVYRQla/JXWyUSwnl+qoZKhBaxgMneQTQNIgVI5FvnEWyemK
5pFpVJLyzv0mBjNjq2ffqMqs16Ypl1fZs8Y5SMfuEnNfbV71slROuxhznXwdtmfwghmJEH5Noj8R
TEORvHBrvTvomwKaj8bUvPCcS5JjWVDlw+zebRPFip3CxaCWrlv5SKEYStGHiK7uKM3IIWDPZKTm
Jo1caNDhEld+xMMxUwSkypS6B/5DnmFSS4w2VQYawkX2R+hqoiLyFmsbuYI28A1R6i5KmSEc2zyk
xearNcqaN3cwVYbc9cTvtQs1LgOeayUqOxQTjqVnNcgB4PnuXh+Nj7PYKDPgmYBSwlu9WQXQz4K3
iXw8HQ34/9GrmACEzsTIVBlzK25Z1XnPMW8mUQDSl61WysIhC7jz5iDDVFBsRgf7sqBWtp08pc55
txP4MzEgNwOYdgNDMRvYKAgVz8hfaqEYEj91W5HFIlnEeF5abImfUnfhfxhku+ePWWp2I3WwG0JN
cO/Eh2uzkAb/wPsF9iSiqsUORLCWmA/KaRFgoHViAgpKW6UdGP24wIEd6fWHzTc0BKWtHlAPVa5A
b3ScOBJRIZ8D5ls0b7X4gEovrqWgMmy62cojrrMXFrbvgQmwuzLJrJiULDiKua4tGywqnF3g2U3W
/5X5E4FcWEuB4OVyi3cBfvE1D2gdYKo1fk6jJQyO81z3OaogsFKPHnvn6WQds6nSeWcaPuifx9az
kk/kJMz/SUpYtYQDTBKNVCbu1b59qBHadOnr8lYP4uRfW9HnP7Jk9+r8BNq5pl40p3yX9Q5cJDys
8B4Bb97P8qlal25pjkA20iABAnWs9KElNNiukVaC2lAdb1ZK3HfJ1uvdq6aDaOp87RybVQaW8xvJ
OPvBI0gfp0M6v6GgyFRTUtcaLR+AZ9W4ZyEigzfZfBk5feJQ1rwJo1hFEw7ILR5OxXuDMRaFKIYk
NcDfoCKSfmGuIxRf1Aca802LfiRRehomwD7PEN2JvAIya+740CvYHkyXCk92pCMrH76vNB8l9vM1
GkUt8+gRWUTIwRMg8pwrPCcFsKPjEUWgWsLuehn9nLST6mkeklFmOXPDC2NP49fu5IB+nzMraZM1
IlxBk0ZsxlratZ/OkiHscOgN3a4+RfvmicmoqCct5fG0jzEGIaIPvTdAwHR4acyr9SAEhTYxDUos
IpqW1buZM8Hj9qrQ87Ax9uDg/4pPaBMYHYb9Fo30XTjOLpC2QDE+9DDX1nrDZxZGYTGPLZBB+l0v
EbKSK2I8PUX5hm5riKV7z+WssK8mIHY0DhIfpYZ17XSARPEm3KOqNsL9iV3zXXr3QJHrv9XHi87D
Ks0d5oJ/8h8lW4YyVJVWZ0TlQYD5c7XLSEHR7XYo2dd1np5GNhRjATWOvu4/FiBJZbn3vNBQahfJ
D7pw99VRDFf0mE0xD+OvX31j6rhgT9MC3V5oi8pts6JyJfvfZeMIMkeo9lwUp6aF5mg5KNbvR2pw
gjWDfMMtCbRPhHZt7NwK+ChJVhh0mH+pIom8n6KXevJhZCfyHpFByAFu9NR/Ik+zbZSsdTHJRRyE
5GNay4OO4PKYj34CHI21n2oBbhQxodmypGIRNAlLPqw/x/do8tcroZV+wGIPEKOxwTAfMD5aID28
AKBqPtUZL4i+cY1t5295i+FDOwVayIU1+X7mY206u6H0qy4CmqyufTsomLL8a1Zf+CF95CV00GAH
2Itq8XisEwiPL2S2tatZwXzW4OcM3ZRYd/oYeWJMdyh8LiYD8luJZgupl6bF6oxz0eDrEN6j8zdF
mHJ9UsbDxASvrE+JXQubCiKi1t9Etf/XOGx8zCglip24zpFwGtm3Rs9p+aL1E1Q9uIoe8BNMUWX6
Xv6xSIV1Do8Qtpvrs+wzqkOjF2tI3s4IdgAEgqWfBaDjKsTsieZaHaWo67oiwtDLjwpKzxBgG056
ixaajSUQ9oTtuID7xr5YJqThBxVFMk397HGyckAD6GYN6nafOYjDPj5UgKBI+0BtUCVl1DRaXBSb
+cc5bcvzEuyNCtHeKJCSpRAaAVoreaRDXuafvYOIBMf9VE6lPbf0SmMcX2G/k3WIFLrbm+56GPNh
r60esoYzybIOVeJoCuOxxtM0qsNI0EOldOn97aQLIwpFp9pa1oHAoCbJqD8z2gnFUEJuS0mwZGaG
p2U8/Q/xDru3sPp69c7AiND/Lnp7UVvgGaMOKuB6YCTixXf8fBcEE/oUNWXGVd6of+mhlh1i7GFG
9yj91dBvPtqZ6zL85YNpss7vIiroCy9A1Xa4IB4WrDtBLINFpJnMAEiN/MB/4nNbSlFHHVxnF7Pq
q1TLy57HDzGJsHQLxbYkgZ31ywK5f4iMDh0BnnDnkWChz/Pv96OdpECm5ZdLvznD56h8O5LCDzEq
Mbpp7KGxFnWa6OfmLPTupD17h8bfVab3PJ/1YTQ2UWychCT3cLhEPdXt04Wb1t4Z0t4mlrDQdQeZ
Ht4IS5SagCa93+Nus0IWlJucrxXvhfx2STwcPQus60eHpXj09pbN52bDzRBsbXSdr4KPkP4qIH91
5B8K+iVD3HL7+DKcvD51c93u7E8jKFPwd52PKWldPdcUYi5ynd/O8+l/EpLw96h5P1kr+Al2bxal
yNtgoDAZmlQaG4lzSnm1dBDdBvSD8TeLQykOdmI42wCbUr4+NLImHiELNyFHIy5tHCs+3kcLs0Yl
i8Ls1ixjJECX8zP+K5HTBPKoA1deJNEPqfzRcvwPLpkX8AZ+BQx4wKntl1N3SKC3QXy06qmvsLpn
rTg0b+li8jvkNgT5fx4B7rDQtq+A72u1/yGUpAHA+F+9+R/pRF+K6Vbmvy/e3cBqXdc3kiHVBIgv
+RhhIBxgIm7C0qTcVPv3vJT28XPgSBRnJRkKVxugoyt/II4Qak0AARn4KrIOKOdNy3YokSJ1PkPl
L5Im1CjjSyQJNLhmqPGZvK3eetPL3OylYlxjBl6l3SFc56lgjAzKl+k1R+QJwtHeq4afVENBKHyZ
j7euG5gd+fWtrbNTS13qq6DTpkQRiNnhfbTWV9/qhm9EtnMeItsMGc6fXeav9w8YRTor2yx4/hZw
RwVCm3sWVbRZS4t/C3hwawJrU7p7AteF5MiMEP90MdEYhTMVBgHz441+4pj6c5eRaO3Izic8m8OK
xnXlroxCRrWh2ILUlBErtTf/u9wp2MBvg9QN7VitPOT9LoVSdf0T0QGUG9lIY+v6n+XuYxGwW/Da
BYA5vvmnZs/sEx76A7v2GiyNofGVXl594LFaZBWu3xUg28rRdrRxd9ZjlrFf70pjlhZNCe07e6eA
uyejmQxm5FZMGS9TAP0BdpV19FIgUgTDTJtaZY0VA8/mCs/RtKHCzi7esHRQaKk7PpGKL5pxwaRQ
GjDPYrW5S/I+ZqbStRpEs5vfbw1e3RWQZVJv9DXfvsiAqO9NADM4jwP2OPOKfAykgXk5VCClMS0q
tBr6b0jPFAwj8BMrdoBzJiMZjvfHofUYWzovGOO8ZlN0CsbT3UvgMM3M7dm136BpN9y1dAAJLdkl
a2bbHpOWW2zpTBuxXclr0HAKcvYmLV6K+5KIEkWgFRgdXAyitXHS9bgRDpSV3KFwo2fkpxTRGVkD
ZnRSThCvFyX2qMbRgZbauFUKQMAlTlyA5w55534EVDE0OSqIh/DeuaVdcNLQBr9Bk+BOGy9KCwPx
qD9rbFqDwE8HXPJ5EIhEFCiTYzzhvDjgfWO2gxS9Lsvr4m73oT/5XLQoubP3zDRJaofHzPTffB0N
tUpKFpLmIfIGiMVFhGiP3XCj2lAetYESMdlwefa4hgTe/j1eSnucKnMSAbAqeFyKFHIVNigq4SoB
NV7uF9UnEOduxcKF1QYw06Ii7Ug/nXEJF8xy9gmLp5yoJr42N/401MiCUjDJDa8Ya7xbBq3RgDyx
2XSXe5L/y9icc6wR9iHHccQp6bjaC4+UhS0yEUVO9vOE4XSoP/Flf1eFbaSRFGvni8V6QvYvJaYG
jn4jpvU8gRlSgjRExGa//nME7Wa3KIU/YhMkvqQI7hprgYhk1vx6RhvstDctk6wWMVxBACdHNO6y
tEdHPGN3Zk+0tb3M3xApFkzY8DQeDcDRD1wQyARsX1/CxrSXR+jmqgfdUoz5yhbIsKTRGuztFE4A
uih3w5hfSt+qiGB7kdr/2ixkrnsVZjcn+LxdXrA0sgoGQTIMr7dRgrPXbCbpuOk8/WBBBA6AIluU
yJ5PEtIGMjKmYjC7Gz2gdT1G/dXuDD6Aybs0VMA1u7aJokMQDHCbo+EJKIIco1KfRbldSklkNw1l
GbA8BQemYXXpY8ck79VbWS2GL33uKG41X5TO+/v1TmvNFDvJidUyjLqUc+3Zh68r2ixzAd74pzFS
Jk+cA4qZA6qPHxL0FKb1BMP3y02q4m1s8p8lFqUb9+CdM6SGi91GGLswhS8U+2yw0XMrf+AgNP+/
sJxr5UXu2Y0w93HPSKxNYS2LSWH4CeGvhBM4kLvAtQKhrsz/S9ILnpNx2v0SlsZwsrHa3hAS90c5
9kZpEO6UiQKckePnEOSgDvrngruV8T2HXAxvZ1SOQmE33cqRbzwFwx5vNxqnuekRJ4D8AHSQeDZr
DV1KaxlHnnD6UiLakhn9BUsqHzS3jLOG3TyKTceO+AiL55SxG5SIpQGeOJGQr2M4JUHrbE5VsXLu
+Z3jHbHxSZn1Zw2p8NU9ZPF8z/9j4TmI9A6uAUjxFl2wnhfsmbBPez/dePLkrgYln1LnEv31ZqxE
d+nKwseNNtJ9DQII4Gd2FJGdQzf/DgD3StixXR6PO4FF15AikBKgcJ5Jpl9XqE9Rl5h4qML2UFK1
CptbKXZDswY+MOUtdKWV409zIj4RuDgHYObhdGSBL1esJH4n7ubdVXCqcjO7MT4juCCT7OIEG2r9
tN+fX9qugljy66k1t8pRC3UeRM5cz0LduH6B3G9oXzq8d8+87nhHuDU3sSM5hxG3DPqP1hjR+OGo
29PAcd3bTFCUdbKEAH+g6WYbFBk7qA5vtbAGyB+fXLidue2u1k6QEeIdnoIcKqYn1mdg5z9ZUsMW
xqQ1AeDDkbrWL59yVrliYT6sMenYiQBktkXII17UC0EaVxBGJPaph+ChAtzgPRFhE/8KuviPkwkO
kDClhMQ9jB7QKDwyvEiLpMYiC1RWLNF56ljpSHJDkdARIQdrYnEPtQE73DvI80LVQLsYGGvQKUp8
giJ1YOAAvuwdTf3STY3szQ4IGc3DjA/YoEw4eYBui1xn8vNIFYQqIOTuKO7Au95e0dZujpAClGTb
QJF+pcREspgAy9s29zFv474W5lk1YsaTB+oIRoMA6ddJMhc/e1BJ+iPnNCy4VDcJRtjxWqLCcExE
T5KDxSKKpMxullN8cujeD21te9fgXNDvIiKaQEBpJ9ck9YB1NVWZOCj+3MAdWkUnI03YYJDVsiQZ
sdBL5T9kBjAoBLn8jqESt8ug0SKaelgCqfkuLled5AorP6rStjvCvP6r6uqKMLKWHQJeIYzrOmKb
/IUnpGaVpn1cYJNcNwzwDy0kSG5GUzmpVQWWein3IElmCXvoeWqVuEVSm41Jb2Fti/t4pvqZX5dy
rMq3PFQe+1rLLBUjeOlekB00tUIruinRlCz8f/nJyyK/amw1dC8uPy9h7O9+3OLvf+o6NfbHuRka
yx06gQOs/XRJO/ej4c4y6KR311uogy1XidrRHoW8ZZBLg12f+k8H7RPdn0UmqgenyYfli0+pKJ5m
iQ08DmyUykjj6I9M4u8rG5k9OaNQy2zg7h81/9oko4wntBnvtTE7BSuK0x0iw5C16RbrV7P+lubI
3jIYzOxweqXboIKezXeIV+9cLiyk1HU/mzZ4NCLgIbTRc/1zgDrIRl3ZmBF2XNT9Hx2Vxw3vovkP
efww3UGSeVbkE/bw1rtsqgi5UXmHKt9gpjug2f62tnlMztqDeT4hcVESXntRLTHLOOLvUbAyAHU/
cf/nSh6qWFTm/QXnU0WXFXgi9z+y3591SXgitO4tkCkchiaIMUNHJvug/0UrBn44eDxlW+htG2wc
/WWw7SrP+w7omRVxnln3ZFk6p0R5ZZnuKe2jVeiIpVsMX4q9wWtH+E/EOUr/vZyDsIYtyhGx0LfY
dNTt/pFhBrLZUkuSP4NnzYYERu+EvcTJuaWWByfOL4nMto209VH067l0exkxWqr9vNs2hOW2HXT8
hecOEZ9R8PI5grKRiTLJyvI6RgRp2KfGCzYsSORImVIZLjpXxR3YxTjGGeX+fJS1p8fLOz1N/R4H
nPtnlrQ/aEyFtkr195Ls7+22ecYEDIt0LiinnEESXh+uFhFA9hgXSQWgT+CPdZSw4PJZyROZw2b+
7M6RcfYaLuyebd5Z296/Uzn2so2OxDaLfBki8JB8VFkmumJvQMy76/jQBAsxnAZoBWBaEIozWXwM
Y3WJe6PqXwAlR76mSY2wH/AA0/LZIRMv9E00iAQrW2BIzXJdE3J7Jldiah3ZFpKbeNSVEXfa99k9
IVmZGIhkNpA1e54U0PfbbpxaVdSlYtfWuuvg8Q6mfRFStNTU+Yl1Ea2wug3guzMKtB7Z38brVean
u3jMNSLY8MuwMuuKcIAWiklVaFfR/8Vw7+0EJU5uqKBnrNUURZ7WDTs3h8GVZsXGqM1PZP3E1irH
B4bnifF30GFSdbxVCEBCbvyU5/7IDazbR26aYWwzgpc9CpJtMzknk9do0pr9fNf2YrRT9AUrGTXS
69PCR/W88vmqX7GIf7DjtNmWuyx0IqI2Lzx7JPZHqRfBigsF4P4ZwM82eHjKd+iZmRBJ2cr5DF0s
68FseVYBM4MKrmte3ft8Z4GV8C1PiVkzgYDd7rIsWoUsSDBzPKwF5I8H5sYKGmEDmiNaEZa8LZPP
YGzLZqBLMV0a39DftmYWMsBgLbbgcwEI780MnvFBfIyrFQ+XQILV2aOvGte7Lr+YmpyK+KKzOgoj
3XCuB87v/4h/MaqShh2wOKWR0LxueX5I8Clbf4JMa8X6Q03OV/buvGhzF6jZLv6N62YnVXoq8tyS
YwZp+OUHCdpkKDmJvCNGMgFN2+dths4INjgBVglqM5OBUG2a92vDpPABOtvzbNeBqxvaxd0OSZUg
PxTUUqyo0FNZX7m1quwpAKYW3wBXshCSype3eklEPQchIYb4uOFdXeJ1a/cJZy73n3FjMPEZvSzQ
pIOErxjeyEajB7WBtPzMwOqoo0Tw3CVgIY1B4xa2gFtbwMRZzM1On6B0FgiMKkb6KQyxMNbexDm/
4832nL4P7Wz2A9Q2KlvoABONBD9UGj7IRY7cjgWplYFLt9QF4hRmdS8bK6bKCOJ6mUTHoITEqMNY
kOt8T2UEwBOG8ihhIw0/FvgfCZSsgqR7wGldlVGJoUzTYwbTxRJ26raV4bMzTcy5ryhEkq2QRJCT
BkE6RoMiQUN2aUXZmmE5897MV46hMpTA6jIMxHbS+uTiqnlduuvhIozXrFVEFOYiSjCX1/oNO6Bn
EvTfNv9l+7bv8JOmRxEBf7GMRVLgsumGgmsr5HFfmC1hL+ITgW7oYG+yodtQr9jiVBUTLu941V3K
JVAJMVhXnjJ9j8F8k9QRzvbnMhzSHae0Fp6sZncFAMQ9s5WfSb3txx8q1oWqpxZUki5YkvaMv7UY
1nQOKonF56uzhwRS/tXrfve1HaKcJksHGo9z3gL//pLoO/xZq/PEfa9eH/3XvBI/LRyFFQiVZmlA
3/lB+veomxHoP592lp36YZijm/9a27skGbY3lv0QghUZ+zXMW3p1IsT2BmQzqWa5ymYIUEk9274V
jiuZeDlQeDxjW0zRkOoBVwn0Yr8Cq7kpc9orG8JyR+6JXHizeGnvoCmS29FwcVmGnLvXrg187g4F
old4BO+MBuwZ4JlR8NO9pcpftaPAWS3icdFsa7Uy+QvUOLv1tTujoEPa90YpbDuixcTUhzwSOyFJ
qcmBkzK4XoA2GAHzW4JBJWZ+4qXKF4MzvLcw7uojw1RkpkvhEXViF08UuD18pDqpgLrrQVQX1UfN
xcURAw6V/3iS4XObRPDbCsrYYII7lyOrJGhlr/3AoNCrdD9IhSZJsFuHrrlvgjlG33TfcFgbA/5J
ZWUBdziI9r93dKhNRS05pl1bxy2skyYpFdJ8MYW0oB5JN7ozOTJpYSchwdeKGFSGXR9MqPl7IOrW
LwME9+mzbQfg23TjJBOF2KceOxxjgnzEPjvKx/OGTpWg5PxAMITCIjah9BkyvTaS+z1klbcavKx2
IPW/4qfgWd7w1d2puejdeFzp85K0nEA9FWZ3h1p52JxB6VdCIN3iIg9aG9UNOvBTnO2w7Q4I10mP
WWtS9wXAiPKgTIyB/nE2eUZvTmAwv8SQqHBWwNf5tBjKJDEn+B+XNMCqpAKvUd1Noc9XrBxcpLlI
h7vx8VZ33nFZhMzKwH45/NaQE8VuFHhsU0RaMKA260ebd30uxu/ckerDR7SCVzynFSsx4n9t3ObR
ruLwAM26cIyuCTuO3QjOBHz02xL+O44ojWIpw3f4Z2keY7NdrDhis9xxg4w=
`pragma protect end_protected
