// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
IZ+jhtr0+LZDl+9/kyD7wNhnAwmYYsdEpHg0/GrNLBZDKkS40JOGMqDSbzAG3sazV8JP+sgXdjLm
IXk/IlXJvNKQMVIJZ7Gj5VyhdpG2Pcg1WU1tgKs+m6yH4/gVh/P1GsCX8CFvaXodhjLM1HlRXehT
wAHjRY0Qwn64N47A4pZGOkGJfYRbmBT/1bXFkig8QMttHtQY8L17dbCm97IE06QZk+28Sp/7fw1b
T0YdlzOu2LMuEkVYXy5msfLubPv57PMddyjMEpI6LAysKQYNwYBgbjHtIyjpxhWNp9OjAsO+Hnqi
CAiPYsbh85uo/UWB0KyjEZ3PRc1v8vsozGlAmg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
Ja0Imka6PwP5W9nWK5ANEl6lKSKIaIhehtyO5pqufL8w95X5Z5ZMj+DJdn4nmEJQKg+rtOM8G/XC
zxsxY10oGTNjuN5Zkg1OEb+4FS+5O6+xWDI40GgbQzHBTZRq68/qvo9nLynWyFkeKk7veYdwgqIz
E1GinzTUa+fKdAh7onVih6CFoiKsANb+1pux2isK1C0/KYSRUbDEdSBENEaunVzltehaqzIvE1UM
W/Nzr5ipWXxyS6TIcp1XwdUL0mFW5gE8q1sxn25A4508nm9awKfkSxfQO6xsYu/Dyp0LCd4rpQaw
KisTWlcB1lthIa/kOLNPWvmRd+6ceeX/zVc5yeZFT1PLdgcETvxtOuAiNnVRJbBII7SWv1jwEb4K
CfcG6OkCgE9Y6YzpkY2+KoJ7vAd7TYtbZkYLlbQjBaYIhgBfgx/y2vIxWqkhVXIaMxXFDPIaLje6
mCKhoLVYwnkhRtxXHAumX3bggjFCvk1cDQ6i4SVy0TLU8wfGWGAgWTwOwEEjNdgC00r9FVstSO1x
PbTYZLuvTu39deyHmVtGq5dM/sDduLADE8qYi9gi6BzwBfWaNy8pClYe699uXE2hNIFwDGZhSeD7
l8dYR1iNta3GLUFBJiwKlPUMRFdiK2/b1RES74f27tpgzbblf/zeHkO6kHzIbPD837qCQhR2Fcvd
+6s++NK1R+CLXtBfozGa5tneNDb+0/ULrKBLqpjRo/JnnnhpLAxfkg+oiGejWtqhOAbhKHJsBCir
+LeDZDBIkWY+83G+or1VtAfPp/uVp7Sn4X2ez073HXSL1ACa/OXmrAumMfPKxusv9eX30Q/ByJ5t
+6WUzbDBsDurDDcCSrg1H2kfCRNsoaBz2+wupIppZMND+mubW2bfbAmsyeZVBSNoktui0UIR5jIp
X1TEgsU3hmnXPnHngPBDK5xLLAjWoohdaztPHrRbR2lWqGBYvAxcfWH5vIwHaxV9BBJCVa9xCXFR
b9yvXqM2JIs+HI+TL5JkPWZMEE9Ak/hJulwIyEModheGS6WumXnZOgkF0vkbNe41LsOs4xt/EwO6
S2KfzDgkM7XntDy37dbJze2cAvGDzjLF3qmhTvd2hH4Z09aKdgj4wAx6P7Tkx3oR5uCNfYKYCjKJ
9LmdnLX+pXqiAnGgvOGaA9kdCqUlq3GHu1A30pJxCvRigqwUkpGbZZAubunrn75gLfGFXR0uhYPB
p9zfLdbYj4Y37eB1D5nkbQ8Q8KhJ8U9eCAeJasx4rRm2SFGWb+ghrsPoKFa+C/o2u+XvmYJT/+BH
ZifnlStgtGbznHv3fjPjtYBtjUseoe9S1zdbO78jGIDqvhBPNRM8FPcb8p78fvbhKsd9cDELHvXk
cQvHUFJvfqf2CoCbm3cSjt524QfAT2fuyFXIulybJeTu42Dh/+EYHQVDA7f9Gyk+xW+abBoGxseO
qGTICKxnA/T7Z8Pn2KA6hAJw2JKgr51c0nSNB9L1lrJpyr3ZMXDCslYrksDJ2aUwfaw2YxklbM4N
iiuwG5VllW4R0eKS+MUvTrOYheYto5vzJmJ5KSyJrs//bCel6N4X594rxYBZ9BhgKgfZlthCwC7h
EQZdNe1UqwdSoI/YW4/v923IQjHpsjIrd7MtLc3ktsh9SxmfTmEdM0r8TaAw9w0xvL373tfktPkR
8c0XylXMDzfmI0yg/1GxalvUasdKhT9EHKT/rw19V7RHFQ7r6oSzpBjkVGptiD5uuR0xlbbVI09V
eUOKTnXgmPYZKjX9SBo8kbi4Mma+cRUCR+2gVK3L5p8QU0tNVLCndKm5WC+P0GwaFRyAX6wfyA1J
im6W9WUnO6wnAM+GFygYptnj3QhIngebVlGepF0PsZPLbu0ReY3ulqfZ7/9bFOJ6eO38f7PLtuxj
+NXfQRIeFK0xR/Nt1tf1Has7wkVPEOytb7TitO59JE9LgqHfI7XdzW7P3YnT91fHbu5V2ETN8yqL
n6/8Fh+Sh9qHi2n3As1fHBaI9vdMuqgOyDTgElLgGuilBoX+onkp1G5MMg7+5ds+g6fr7qf7sQDU
B0o+B5aYJsoUADLf7jpzXqZwvX/3Jo6UK+WayEnEQXNUeFF+i/pBiZSy4u4tJfVoP3NKKgGCFQrl
laJakUljZfuqfaMKSZ4dwaZoUiCpXT7fh9KKFCS6PWmoMDyaic3O2eJhTBoUaMf/N6H5Lv6vonVS
8bbNbYIpQGi9xpILT5kxcY7kJQZGjcMSk1l0K5hLeXaTpJGMNvqrN8iwz3A0+7fRw/EqVla4wPLk
6G0qt24RMH7MRz1Jqe5ypY7tl61ggmOCEBl4kN9ibxD4jD+TkZQZq+fZ5rM9KF8pUUoqtkacUuYA
Xv+nrfFR0N6kYQGLmY7yED38anyt5787ByRth4LBN+8T6apJNr0Hp9C/MM/1Za9a5+Xp1moMLnIV
G2MadD91tJsDYzMrahF/nV+V94Q0MoikNqUkgGsNTLot7ZjkThSfSng4IJg84n1vQUdNEClVqX8y
SnzN5yOYwtxv2LwdFVy/9MZ2QGwtyH6NNTprXFCUQyg7HyU2pi3mfBcfC4AlZm5KRCfCurx9ko5L
usmd22x4EuSjqU0bwLTDADwF6q2EDgZJIAocu69N6r1lVA1/5NN+kTXRAR/IPCWcXzWTX+Lf5ynK
IvWDczZBByJXPPfx98V8NbfuzcmWHAXkIB5OYmkG3wwNfMRGNeTR31qp4nr9saxp1C0m6RsOEoH4
cAFytxb9bJHpNNYDbeKLjk2OjPdnwCAfGu5lSkTkKoxNNvf/vWPqz6rtpNjKU00EyRIQUOgNT5TM
W1h65R6DlibrJE3THCLiH1jNPv8YqvRf/yb06fc20HSqrkkp84V1WyyWPCKmnLNYdEk60yAf4TBa
CU8ZoQP2Fwg2saOztN7YE2kxsvmBahhoO+LSaVzUiuit3p41uh3PMsV8OnkImqH1R22v298UOSDS
F+ip34qgaNaBCs61Lq+ZPV3qQfPpCLMhgp+VQJnEbBHHKzhkCM+LaMnU3PaqtrZ2jM4msvds/oXl
epDkU2bfCI38fo8ab4eeJHRqlMmy9pruOCZlJPp3polbAfZhpDkOd719NI4VkBdtV0OMe2lGs7Ar
157gFFx1DU03G1L2qVBbsdFrJTW6lxMlxCUBLf82pYVGTVQyX6i5Wd9fbhUGgJ85D2+tGUiMQn3D
V9nkfLK+r80SmthMlVqcuVvfpxD0NI23UDTmg6jgmhV+r0ygaHiJ7kvO6wNyEnKKzsOR9QpA3ZSy
6cglNjlw7xWImlC6eAnXunCBabZCZJAf4w1HIjbOMm6yQmBDIxaO3wJ9DoTJD/QV9XBDSzcqlxoR
fSAdkc9w8phJpzy7tuQuMj72gHe35d/MQ3bBQNwOzdt7IwWD0Igj3Ap1YcP+6QFa5ktNle5cRmyG
YD0mz8JccoSWKRTvIhsnQBBZPpEG0ynhVuIJmoQ6M+EMJIP0pxKSO1M7ctiCmrgtbMH8RRpCce/i
b/T9hse0Exg8kcoZxvMytPsB9sHOmPbnDGzVbQIb05yZlyYi8pH5eVDl34a9+09E0y+iYSo96KOl
x8xU4yTHbh0SPgiwUliPNqWUu/1bqPbpcVREZbi1v5+y2VIv2v/ATt1N/T+RoFHqHr/R3HUqSqOP
wk7FZo23/8U/StL4SaJNegd0uCCPjZoNI+y6Q5Cv//qbe7cGCh4gjJtvsB0zZTqnUE96vgRrSNzd
PGMpjkFGI30NpW1J5a0bbLM+qjhb9qo7HhQ5FjO94Xg2ErgdshIVF9yGqll8xRyIrsV9pgoJVqA6
r39UxZ8M+PPtL2J+G6rRhodulAgmYNuF1PeXZHRyEtfqPoAf9do87/LC3J4bsMIJqX2APcphZPAt
oZKDTwFXVo3gUTT268zKA4BdByHcohbzusaQwz+RpSgJHasl51T5pZYmLa4HxRlZY4jaJekirV6N
z3MaUg+B/+RE2zqP/PJzXMGR82bNwYVBKq/X/hkcvDm7epk7Yg/bih0Ix4fHpBW6oFi9Khk9iRuD
fDqdRW4ovwAcMwCSjDWePA5x1pSKjv2qlwdWX80JJ93ZIt+Heu1KuTfDvqd+EvAI8QWNMWhwSfgf
emb+a4UGH8M+V9dm5LcF2ZB8Mr/59Axg+VhySsAtd+UMnEtKeAiCZyp61PWoC2QLJzGhIQdnBCUP
7x/zEiZQJq55DT4FsOIqfiM2+wZJDfSvrYJ3OKJ0VfkLgVRd/MvX6ehwNCkT9kQt1HguJ4iwhMwp
IwpdGkJbx8HchVk7LkmjbW7qWdN5ykhFkNZV0QTRJJTDfYt1vIfG1dp7EBf16k/oRWS7OtQyt8Gl
7OSntL6CqymFvO5YeIanyj3e0VmsiKsZDde6x3wnWuqVRKX9rTa4hQqlP3mHTcQt55XG2KTABBhG
7zrRbUiuDMOQIBGAcyVNUAxOs9whZCs6NhhMuwcZ9kJSb73mSeCiE07MmfSgwDtCgBOsgtBUv1Rc
/zyKWvoQ3vDSrA7n+Wm0LjNiok3eqPqPLuZk1jpxnoKqph/PkVURkd0xu7niySDO43l5c5t33+Ms
0djIFdfmIfrCUfRZyFWhNcf+GqGaY4UBZWWdMFrbqRb6mGpyzEntPhnOPZLr/zI4fV1VbMsaHckC
NZyQlX7hbVy6QdiH0j+BQQiV++MjAJ0ccUNDUQrjDTfV5mpYu7unytLgFpZo9J25tmiXW68bol34
mHyg5Z1nGDDtucwLMPRrDHEJ/3CH7Qe6k1gEkAwPd+5vQU51P+wykQrOHW4VaozHyO3alzPDWHic
kjF2Kty4jdOJzG/VCYM6u8h1tkAdqsBwcJeKr3VkGC0DmMe7A+lXkIYscXbxd6J7sfMpQvOtuUb7
vF+exsFKKxWhbZ7DA/NJtKFuQYlNAqpwRxGwWGsY8DaQa0O0Wy2QHaXCMd+sJNnkb1revYiNrZfx
OckiUu6Pc3js+yS8CJ00GSKPgDrsU53k1JE6vB8q/xCOlC2k1ikT48hb7II+MrO+y5J16Dqcimqw
lISfDyTI7rImedOhDinGXMcyTfMQBpKG8Zu87/u+Y8P10n0FCwrkeie+mJMME9sUZ9GOqu1r32X/
uueYFWxAGzvam8yrsa8wTfKg39L9uEHPlMI3ukZ89Li7ZWudMQQG7J7ccbWSNDBkaIRs3KIP9F9s
52m1iNJ6EHZSUKvdx70RCHidEFg0IZOnDB36qPTSIwCtHTZhRhrlaYj+qyyOqhaSOy4UPIBSZUFQ
t6xiYk+0Q1uJh6mxoHvRzEknj4+CPDzt1dWfTcsNjErSFedKiEBh0kErkKg4WA0YsRJySTXLTpYb
rd4Xg21c2tj4J/iXPIdUW3RLWL3z6VkdDBweHIBOVuwe9qhdppDTj8apqRgPVqA1Qsy85xiwCuZZ
j/h/MFAx8Wvw7xZcQqins9u1A+LgT7kRjmiDiRdr4Wt7gIZRB8KgC6nRB55+8M0/if/GglE7oSps
fe2XE0/mux1wvp/jl/k1Zt00IhCX+DEa9Vrs0lFg8iiGuZCyKTj3NyznVCNA2hjkN49t7Ie4i9EU
Sdl7wXWypDqWaBCzge9GFvXMwuih8wize17a0cauBXRwDegYnR9EziPE7ZaHmrfJYvx2iGPD2YfJ
980nd1gd+qp39ogjxQ0fbz2xN/2iHrKmk6miJ481bSRK03qIJU5q0ndmJfCUjqyIdpe6sn6akoeM
ZFNODbkhOecPgnhBkG59VkMY5jpndEq+OoEtQGbFHPCP8VMDSuQnCLxIRaQn972bSsePIs2R21DL
nZtWh7e0+Fi2l+Ahl1bYnF5815frvsU6BlZieAXUqJOu20Fi2sgzTrVY/JQgsg9irFtDH3eldGLO
FyxN6Cua/86rI+5tySgtu8udCyfDYce5RU7elI5wkeFhzE9YJIOtMv7MhiOFX2uB28zVqZvzhCJq
9lY8EmOkQ/I1humKTmYQm7QnPXhJDOdxZ023l56oQdD4zlrCqlUzNPDOLTEYeWo/Xdf9+nd6QNG+
9ELPexX3T8lEKkAoXNiTefOQp8I94MG12k01InYlwwAvzlt9iQYCYLxzLBkAwZiVMeTnvq500tDM
rig2CwVN4h3Hf2QbwKTDt2nW3tAaHKzERVhelKMISIOJoubdh+iCz2ox3zcHiGSxJu5k3Kyhyc9D
UbdWRulgBLAekR7IzVDgwqNoJjM1dSwQe3PM8egM1lsPY+Cozuetf/K/DV93efv8d4pum9XdORSj
nMMqmMnU0LR7OcDaDb2Rt7AmU5MzOTgKSzHjiCUlOEzuFVUt+VBT+a19B76qZ6Y4/yEH3b1WVck1
yyGGzVF0+zviRWFXBprHVNSvuqxriJr4NKweGnReLhR4bjf++645t5JiVn1e2q1gSz6MhQB6OYv+
47eX3n5NBan1Hw1hknnxj73AoOZEgwMhXqbYSy2HeYLfFeV63tucfj+VA8kMSRB+kjUE31ztGztu
0XdDwq5HI2bpMRwd/heEst7bUimOURd1ZWWYHj0yXcjn34NImybaAqSY2Q/HooQHfEN28fu73ZYK
qv5LuxQIprj5OMW7onPjjdgyr2hrGDKNOxuUQ1dzOmFEye0qM1GIaqYms0hW/aDHRGiQ+PGaLeSc
5Jdcu4GS8YbeA8AoiSdVrmNcaSnw32FtbLKvNlPDSkLPK4zT6xmUY0TSY/cziBCT1FNOQhRvMTxY
T5mQm+7cjx+UGf2eEGtTFBkCqh6R4rxkSUU/QojVLmNXLLGw9lGAlWKu4wEcQuMY5tKOV25yWdxy
gd+VcGcTE/mZ0SYNflfONLVO5BfySYi1mrqZrbqvVyShzr8fqwFy16GQ850ZTqG0p1ZqocPPpnVY
7D/hss4vdbe/coSAUbQ7JzgWGN/tTpJuFGcsGEcSggvg0Uwy9Vs3pzMlSwpN/0lp4gys4ekSzpmy
86ZHwE0JpFxrug/ap5BdTgKbxUZF6PuygZ4AhuRxcvf0/LYDqo19AvAmj8hLTxu8DJ86bj152VIc
u7qFAtQrINFibgoJBfzK9v7aVdZ2CdxvyTreRYJaszdQSc4YBw9VJe9+HC/rcIiw68d7h22vqPnG
g+8+Pz1wAg9Rf+dA+LRCgrjhDueMxvPwA2gCdvWivBahJXR0dfwYFEhYX2twVPPEjAE4OoNqkDSz
ab5MMMo3PjYrvBm1VN9j5+QFbeB7padVBYcdTw5DIJFHSdhRQRJb1LW0d1q39LY6tWCMid5E+5s3
BysoQRdwDiucTo3W4vNPqXpwDNdpKTN7nzEqJgjN7UYgzqXZwMGLW9rFF0rzrvWJSyfOZTcqB1cM
qPF+LvBKwR3YcvobB81fpD700eBHri81AZs7DZPgR2iezoL7bkVWhRQBMiPdcHVLLtovyexj6gUM
F5+fcJKny1+cP42dA2WhtVZ3rCtgtBAL3heJGjXKKHK8RXY/RkY2Qzf6mZT896We4yu6FpiFRIOu
0x4d1Ug9R+HWE602Ah2ZYrRX+dn500GmrppG6FnUi8OeWzFZ3NavNeTDEpnrEgKR2M3ITXGtUC/d
230wpfU+UvVAHJfkYD3yv5DrLQIV6rHDM1tdgyUyOW062Duqiq1qoO0q5FDSR8WQxre8ywVQrr20
YHZntMt6MvVlDG0P0gNy3RRPEbefY3uluWccyfEvP3jtwlTIjl4Tes9LrDSoSrpz3eF9ApGCBUXv
iOazTWA2qppjy7uHJN6+ylqQDLbTmiviBR1XY0wk52z8I5HTC7qGBcfqOx0b1GekZqa21kkVsx2x
B3frIJQRIzZyb2Dp8xEqa6V81PXLLX4/OvavLCP6SEkOxE9VIWgdkp9ycjx2kWTqZ8+C28GWlLKr
FLZxKXy6xk3OfHoonBHUkszFEC5MZX7mvH0VUpcbiv5WF8ocxYpvieHHY8BhSGiWhpEVOOL53Z6F
xmJoiZNqochBoBa5dCMmIssPQ15Mr6zyt4OB96s04VT1Qh3cJA89z1VvSDuii1YJmUvOv/AN+MQU
/V8lmjB3yigZkJc13TbsP50dWhHkuHXcHFueNDM86yGx0ucUgz8Cy3z64BrHYrvBiR7PQbDeXXz9
WmQTXfORydMTXdym7WopsU1tBB4Gd8kjxkzXrJkVsn4bvV9fCZ9fmxCeJ3ex4KAZrgkSpfnGiJ70
Lx+dN8NpD9fiAUnAVW2hi9YUBJaRIXZHhC0EVdR5g56BZF68s0ZGFw3m7bsyUr2yf7Z+9gIWMLfV
5zqVJIxGT5XrF+TkiLYJytb2TAX8lTH9xTUbZFAGvt7uJT2S/uFv8vh4J8wioHGvN4K2e48Cu27R
gNUnpy/mO72G5TrUSyvTTDz+gKnH4+iaQa+fMCJGhSPPYY5X+bHK9Z+Rlb+jat+xNxC/vp8XoCok
BjzHPcShsbCA/q0vfCVqZ/qu+7rmOXyqDfJmqjB0cZn5Tap7iseWMAfhRdzcXnaN3XVxOiqshRZw
zNJoPHmJxfAN3MlBmCCcT6AzvBMujF42QLxMHUDXFdsS5tfjQJ9zLLUyHxfvlALFJDpfZWWMY+sk
mPx8g+gzircgV5AHFBa229/M9OC1BsiyqtGe2S6MzbWpEMUPr46JLLIpQ3SSgPN4WMaglJgbrCJj
H50ETDeb884Cxmqz5E7/yTh5ROYS2eLpl1GFTd2vHT+ZwkQCKO/VfK68KfVxc50AARnnwZOu5JOY
3W+AdSFFhuFm9d87j19SbC28rhju9KZxrN0rBvfDh1Cr9T0BXdM2KhALcu5WpmY9X9kMs3yeoadA
xj0BiDUsX7In75vPmSk6IFuz/kaQfjTvIk8W3XAc1K4+1NuYHogLiXy12hZAeZ8oHZHjq4O2/Pea
Mzwl6q2BkI+4jQNiDsttX8YcSuiOKLocQUPIUrcXdckNcfwxoZfyO5kUeCkztp0cTWQtdIvOElGB
BfiSfp/DXXsQ0RCJ6d721UvgfFAv9N2O7UnzDR3327SDokPDtRwbULzl1SNeDpzbUJc+Clsk1DJp
Ck+KXiwnmm73cF/JEzrlCkhe5rRpEI75n6VQmDgSwbk6RqztZHrtq2a9SUu9ks7/DqcEfzx1GiBA
GTWdkgFHLMLWMwunoZ4XCEjExPxPph6LNPejB6jCwEmNWOIQLMuf6JHE7mP3Mt23/YrQjsQ0etzX
yClVjr7UKhw67F5LRQAI9nwbBZ7Yu8JgYxkzgs+mvK6ySMi4Vi0dbyNBxCI9nhYKBEmUWLccbGpy
KUH7RjTdtzUSZXSSAPfN/we32hYqj0JAg9TLVWliXB8k6QaZ9ZcTiP3Ltkf+fafMpMZniNMrTKE3
x8b4svxcn39WVvpNg9eetVaVBPgUZMPNwixP/moam+0+RVGZxhJWjlYCq65/wpEf67/SPROJfA1x
UG1rzQZ6NtRO59PSvyLuT/uIvYyR5vvoiuczNZ4F3HLui0ljyJhsE1RhNRVHgnH7Dm/ondeF/+l9
9XmRVEbKQ9p4S8+P2vJG20oXuU9xAvWt5EZIdg8JwGQkCSry9m53mnaS0Bl3mJ12G4Wf1VdWMdp0
nrxyeL/KGx89fpp1yhvzXoBX/3cQ8aYHEusuOsZF6hSzbWiSsiDTuObosnSNNQd1GsU/pHwwSghR
UdFTfO0ZlgCOMVd4TTuqXEq3R5DuTKrn1nA0Uexqps+YuslGLOM9ZH/4n545qHxL3wdRgoSoGc7e
BwpDB1bEGy7gedanf+hO56BuisGDdaRwOlvxGhQXrExmxcooSV0V8uyhyThqjd5q6S150eRNelhH
rDj/xXlo2tLmT0NWY2wBeqMxfxxMNY4li8epxBTvimL/e6sHRjrsFLIGqHwqNQGV3QA+FoYnKfKG
B92ftQ7UFc94mb3ia+VuJd7AR6Z5td7awKh7upSSPwJcv4QPv7r0Tn7YoLLa3Fa0yOpUyPhHJjN5
RJ10vN6TCn0vXWukhSFDRiYE02tVkvuZtiVLTuldTSZ/AMk4mnrihaX0ggoHJdgx1Akbt+sU3sBj
UWIIqjz1r0myv5RXwenAYRWm51+vYt2QqXfDBSbWmciPNaibw3HgbIIs+tF3JhgFXPRfNdDzPoas
RSQUII8eHYibQouBUGwlTLhvllAxMGDN0VrqY+CznXnVM3XRoNC07HgiH50CoNs54T35CYoC4ma4
8V5xDGl54mkwRZA1amAE3B3csx5uCn5I7AGadZvJFqw3h6eWkjEOXIY6fP7J35FBrt85Jf3qxXqt
964oezibks/4EyRVUczIzwkshDTE0+f5SCrbyrf1wwDlgTijy/lvWJJ43SH1ivGXHOrGdTje60Lk
AD77YfERwAQsB3Kle5iPQ8rUw0XGZHtVLIc3MBAXsP8m0k0pTWrodtHc6/KM72KqPugOZwqo4YgP
2yIlxLjOIEGlcZWJmKdssJI6YNwJy0esDzOwZ1L2+jUfLE5QWn/Xr4LwGvGHqwMhBS/LPfC70rkY
GPP+s6BW9ikSWgzIAT4Y1mBHXV93Fi9VsI0Vw5xb6blDxiY4y/Kfjw6Cbv6jKAhogPiSZnE6ReiR
Dc10YE3tT1+57hP80RO06nweyL03ATT1jC83WXISepGQSGUEhEbetU5vyQKEnFfDrOt9lgKQ9KDI
R6xuevRPHHfGWu1FkXxUSAtihAKewXA5EF4koB3jt12g+bAINaL8m+BXhBMaUdT5Qd3K7MOtgIgN
FnN5ufeeKOSIJZEMkve7XqXzgNMPNpDIP4tFT8Xs+FVQojNwxTMX/i0HuM5nFJZVXdWbgQCY9riH
xEQmLTH0J9Iapmo3k57HxCGF+7FEXLELyneEz66kz7IrustRv9p/TyOne6btuMk094WoFkicbpHv
YAjJcLgGuaBNG46VMtXn0QPspZ89GztdAEVC5VDXZE+JtrQ78B0+MxGEQUSqaCI+bICelAbu5gMY
pm2083kYPaeCFRFJOw6B8Dd/m8WgR7BUqzJ2FlmjAdoNygoXyyvJcoxamlkb2uK8bpbGJ0UhLKTP
E4v1vFx6AqUpMKh08rWRrVQRKfwMiyUh1qE37jJ/u5R3S5luAvJJMxoe4U8SNeUB68cnXGoeuubw
tQxmvin6xvv1+17Zf7hI/D77+Vq348jBOxmzaOiajZZl6wh/YG3eg6gtnmUwxoCnAbTZBPnHKw9U
IyZ9iNISWNmWfEBAN1IpY9SFsGuRoVWDXp2eslrEe/EDJ6NIbQc4x1r7PVOXREjcbEjwtTENU1Gy
7xnC4nA20yH7+Ne2DG9vTdQBeF5xzsv76fg9J2CbuJBerYB0Q8RrvzX6wA0qcpmMjPsfsBRfZZ/1
8m/YL1kKcTm08RqM+cuCLDAWmmwaTEY89vBxnpbbyQf/pCnsLzw0V/6+Dx8K9A/LnKJjYZZYw7+t
Dvs+mg1uqOCESYf6l5I0U957Z74SVbwUFw9Uc/dcsdkZM6O0sYvbKaZRxHbuXazFJUQIjGgL7QkQ
PXzgBqJOkyks2VwjMbwRnwmPM9E+Zzh0YxmFUB69BCj0iZjqxICJn8wAWjjyvVz/NA8vL4BfxKcP
zY0hE2JCpM3J0YdTdtCIysUlq6snSxJ8k/z/MpzUIm8HqZW3zwHH+LjEEepErHGyT6DTfqs0Q5W5
IbMGMzDtNXQdr0Jw4XDaZOOYo5ix72bmQy+aXPn4a969IO676ndWGry14Bu3WzVg/kT4Dp5x1z1o
kwEeTzHOsUX/gPpDME2iE4AKg31mJvSWXqbU1+Kr5MiBl5JPg1CmIDZD0RnExef9FlOYZVNoWSGa
58KwV4EMVsH2FYF+YpiZ920TxhAChErUdSZydQfstQQVxyjfn+xAX/1LE3FjXoLOnTCujxK/9hk0
wrQx78WoANjmIeDe9Yx3tWflz+fQ1rZ3qwfD72tguwD6WIlcUAZxJH6/HW5N60uGxJTDaMtH5SWK
plWe3XXO5l/V8MhUSIMeXU+bJHX1tDocG3J6FZiOrrhKT2eF6pB2f9lfDwdtSGgTfhPlkjZSc3dU
g0h3kgQcYHnwNmclOm2+FzkIqftt8HU0UorFB444YuaeeHjJGOQU4spkSCL0ElyVmuIiuC90pVvi
KY3vfheJR7R3X14DNhmlXCgFO4TdIkAoCoi5fnXKC+7PZ3F4wQ5X/xX3jqeWtIoj3ZtIxo6ecAg9
v6C84Fpj3TX0cOyPtN4be7ZDFvhcuvAtptlsHjk6gMEgJB2fgl+1cSljp40QnyzuvU16MRAnLMIi
B1Z2BmsBYmTWmJz7D1zoWDPRA8VCa3C+fN6J6V4IBCm6d8nA8dgZwIfZN3FNHCs1xc//WlTvnBq/
Wl/CP1dEmsmk9dCRf11oNWso44ZV1tYYUNg7BogeXo1kZuGzACxSjFExuJTPxzqtpqKD1NG7ENDi
3mwH3STqqNExbundRSFX0UY2XdFDsCpPIlmaWti+3+WSsxw3/RmbVU+AGjJLnWPQxW86J0PT8Hxq
DHw9q1tsrzswasK42oU6GqU1Wf+t62Soh1L8Ru2ez/+FvCY/cbd3/Zc4sgaXFZ6uG+GTN8llzzIa
BicHXKwrhjizXUGQqTIvXMCG7eytBvIkHLG6XEwx4bgihf3YJkabxL1Jf3CMvs1ugyj85f+/upPU
Fz6H464ZWKGpcrK6rn03EKyqDc+OWfTQVgJOof89S5ATk3KaxFB9ATO7uq0OUDabrGgeotTX1bF3
2AWXthQMM9tZqQQn2U3r/Zq31z7LDnIH9aL9OIUBEOJ+L+yxEJEtI0az1aymvAjAMksr6KUXkgSU
twFl2UysFXTmDv3Kz0OcimjmdXNZrICXpJa+Zc//tOeiNmKerkEhHFLOCL5u/sj1zRodh8N/8S5w
3nixgBj0G0y32Se0k9nCsjotb26FSXsR+zsy4wL075657hV5GFiHti4RiTwC9tAdrgexagHm5vrz
fPGijFv9ikfX0RtEZ73Y+5f3Y+FWyqG5U9dv74NNln3Sbh3MRaAIagqVrpTWvzc5mbLE44q3VCdi
/M0poWIvIPro0uIxYZgQ0o4iJisY+DoWzzm976/FHC5OrR8C0Ngq/+YOs/qzg9UknVGi9pELsWGH
S3Q0cMuNvlRsUbf3iRGGz5YUc3oM206IJo3tdPG0NMOBnaXsx/oKNvmGT9FKfjv0QjcdzWtlkGY5
635kpyo3dMXjYl7SEPabN3nxLTS3VLsh+f9zUsgbreVRALlAeTSI/qgZb4dFYoYNxfMCyP23kIn4
ZWIJcltdT2xCXUq2YIgj61f1nBB7b3eKy1UgNVpgTOcvOgdrn9BHMpvixzi40//YAlWRUN9LSUcr
kDO3zdTLQ/zHt9X1a8RUz7cood82PEPzYsw9JxNNoWFufIbFoNbCYwJMuFQK4IWdJ+ygqBFEeklP
cEfTaCI3ziXERmdgwofXVmhg1m2WdgSZrLyU5KsNUdGGIPL0wIfirJfgV1U5dULyWEK1UXR2ZkVo
D2ocDii8cWccAtWH25gWNF2J9BO6ljUzPch0UozNAQD+ky8bkSgTd/RqLuRvTbPUdQgeHn2kjnoE
J4ma5TFSApzoHhXsrlpXN3ifOc21pEwf07V+MpVOj//1Fn1y1i/GjbaITu+GUF54t+mGxRg91zWF
UrNc+uu7duzkIQcFBmvZiWsH0zzfGo82jUrpG1VuqDWXlnLL3CwSldMBtJrxZR2XfN5i2OT42j53
yW8I5HFYLWHqOsiwpkIF6fd917sdPl5eq6orURbQTq+cV0CI5Y6Ms9JljpKwOApAs4bNCjEEpJ4H
Z0g4JCLBIVuLZj/8J0AdDWj1MwYlxYYaKcVsBxI8bR3+DMHBshmiTKirDs4SICc6PzeuHPXIE+0T
0d9m2nxvlWMW4vkOTqrOcJS+++eT0ekcknwQTEH9E+eKyptPnPzLymOf4Dek1Dd3X0gffb8JOPgN
yTUyBisTkL+iaOHy7Q8C7A2Pk3WcxRqJ5+vkmFMZ61W05uIemZbc2eWSLW2/k9JOoN1QVDUiCQKJ
nKZxsXhihh8GJ8kECX8h9XuxHzLoMLat/SkoUCHSyaEgWT6JZZfQ7qxhmxFpKktS9TkBlhu2hO1L
4n0TRZmLqbDd9V2//kpIPIPE2KhdZXU3e/7aaiu31mk4uoyGepGjhNN9Vc/LZDbQtdPANAsIXtEX
awm0KHW+zqfMM3fxWbKKs9jhxq6cDVR2GElxWfVM6NWWSiclUwoEMA94Y793sVHL6JKKxqVlwVhF
bFNXG02we4iwsDsGyY1tQ4h6457LSM+X/SF1VPvHmsZzHa+3YF13iOaHHwIvDNuKdWewY/Feitp1
O6howeZi9dldNLYuLENCELJFsUpO8DNF9BiMIAbTQ0iiVmFbkmkYtrdYjreWd8cIPrt4HZwbT39A
gbGF0HQj06/HKmX2Q/UkaV27kK47wY9X/sEvXj9ZkCpB0VbEBIi8Xy1a1uOuitioySxOPHqaJ1qy
UTbEJ/7OOM+w/a7noQWCqtEsvW4UME+4qNAFEg3xZUebiBa/SYJ4ubuCYzp2KftrdUxBA3t51PXN
h6x4y6MmVMnVTALuEcOM/+Xchar3PSxp5YGZyD0+exH/E9U98X/JY5KoIEq0l0ZXAqFo5zyR/l0D
MBTmLYsdM/W9OVQG6wpCbp1vYIHbqJbUx5HMToe8WTSXd0Qy7stv3gpYb9PxB+mRMMxZupG34PmC
IIpThTA+FTgesmhIAm5CxYyeMFxIXJJ/Ub0Ii7sC43gWmnei1xdk+R5J3VWFVvNlY00iwczvM1my
ZiFTf6EqkqTGiJlBgvjDYFxVwkP5sTxLuitjgAAgwbccJerIAQvF6wprD7R611ADdwtq5ijPvdQ/
WWodD9mBt3ZrBzKPafO/jXOC5b+E6xT5Ev3s5pi4wiLipc9v14aYMiew/eLkQKm/FMNYCI4Pd4mx
Lfa+lNM5Q358TVta6omKZ3me7wj4/0gdGrg5KwITI2QdzIqHoYCtHzxjlzvuzhPmsMumTjJNy311
KH5hSTbPO0kijgbkySCX6dPZK8UrBE0jaou0GBauCYt0gZOfTg5qG4vq4ovt7gmerBkDFxRUCHNX
S30+kJMWWdvRYFGfxhMt92BVTkWI3peCWRFyJiVv7a2IbhoCAYET1v4HQTk/UNIHm85rgi0gy5IZ
IyfCE1VejOr5LwHYrh7a+bFHY51J/4XeLK57B3UuJ2l64dqe1IoHNlMX+rbUAA/K6VCcOZL23Fqm
TVXcj3+cfnkcsVbnpT7OLqmWmIolkojcWAJFbYy/Rl7qUN1rx1OqtsxsMW6g/gsenj9iBq4PV1d/
qC3KRCd1TW8j9NI/D8Qviudqq1JxcIFmzEG6pskC8p9PoTjCphoZl3qcu2SVw0zbu2Q5Chpt0Mbp
kZ3Ucwux59DfKVUI/XwCeQQpE949Y51IH++Nj1RTPwnM7co+sgsjn1m8hywrbHkmFX5urTagy5W0
sN7e/YiMOukMX2aC5S6ffjVAHqw4erjR0MZreqII4yflhb5Ef2p8D6CPTYnhausf94Anp2ljmGND
hAy0qj0ySsB0UZWpyWxrzPZffSVCQR2aHndcedsOwxfZmOTHBajCGUmCF5DvTDh+WES3SKVRBUXH
opIslc4I1ss8tGHi9BIT+/MZv69TXeU9d76S6Nk+PvLPfjeHF9jKG7VtAHlOMcI39WV+DlQfzZCU
Xmoh3EryGbNiiJDrmPXpKVq0YcReFxcB/dd4sT+LM04h0OxFZrClzRuRCrDSEq+ayM/uAU/NEQ1f
3E+FO4JanpvIOOfA8tFWik9IkC6FBdxkx2DUD321LCXDS01d9v8dvgHSMSV9YVmKu47R8GjB9xYt
22zjn0EDPpA9t/VTQ2/VUJB24SUvfeR0tKXgU6qc45YCHFHGFDE5IpoVB5d1cG4t3ET369tKIVGR
aiUuFC+hP4DQC7IZ9bpU7+8EttrWuPSQys8egR6ipK+Z0h4RuKmkzKGT+3l5eqyCjBfJLeOWlDOe
6s6oIBGDIex1FrZgvgpvHN5uQVPYZ4hKZ5NN4YmsYVzKaQ6dptB3WaP2JhBuvfX6mnYojiIAcTqS
jyU0J93zr6RBt3SfVsvOzjC6rBjxdPozzQLmY42chZX7aqPccUqYAKiD1Y6aS5aa+wL5qOov+li3
sWJoKWjovYJ5Oni4a7t9eLjn0eTuiXSygKX9PJxc5IDf/i75lzWc17Jdnr1p3ZWwr4NkjgvMhQJL
z4rhEhGZy/m1DUPmUK+scSeL2fby9BhdVMsdBsEC7V506XyVqfM4GdCgudS8u+kfNm9DGsOGRz6E
ROag571BWZurSqO1h328jyDtU0t3Oli3tOkDCcb1tgV1MhTPl4lkAEGrcdmRVe9LY+kAud2zyP2z
u5n2CJi/l3+gg/75rglANwRZFlWgqM0cfV81vzMpFpAT+YD5BAzZPrCpJILra9Ips4u8QYeckXp4
mK2CI8776hrcYM+Vqf3PaRDKWGiyt5/wq15qUa+EK2ptexf4K7muqTjS6yCJU8QIs+nDw0I3NqSo
1lFX6i22ZGPoxdAaCFEd0sD5LDU/Qy2iAoq8gK8bdqicnndBog2U5XVwbfmDP0SJpas6CEf1uuNh
xmuu6R/HlkU++yQNVs+LhdSiTWi2TfmrKDQC8iV9kpjkmipPDG3cID1CC4j15f0JdlomgJAOnuAz
iPKB0Y7pSS/7/jvUltBXTuv/G527zC1AWBL2HYQv1l+MmJu9QqX8d/9RX/LAU1E1NOaen0usiV+H
17yP7wMjl51/yxwTgHJfKgVG1QmWbJZLT461L9tVQ44M/3BRG2SpdG9FWnR6y61qN2fBEaA3x8HC
zq6fWg2YTdCvbzKKcpUPFWVJ99KZVgC6/olKeROJrlQqvs9wOpZlEF6lRu6KG/224z0jJKbmMsHS
JhLLbdJmzUPk7hcBiUkxWYD1bqL5yWJZS2K3AorV2gVy1Dop7OXvopKNnt5TSuRWlh+eTuL47ISo
7JDLcwDHM7HaTBbIFPx2di0Sf2AbZgGsz5bXtg3iC0XjN3vFDsDAuHaiASu4GC6Ytgwk7pcktFc4
RhcfuLRZle7MCaS5C4IeG3NhG9tH2FDJ4IN5moW7TjXTE8ZgpJDEr/Qlrpkec7T9A/LIrLQVPMOz
R8EixUJM3fcBB9IPC862TwhB6HyU1EAJ9tb3OdfyPiqq0xRjoQINNZJ2g7GWPm/dqN5PrmDg7xOK
Mx1pMLPvdYsCsyp3b8vmQ7bkvOvZrMlpxhRpDFPLe5/o9DytqCvkGPHS1xhL6NmZgHyKt2/LmhXM
vqyYJIxKnd61R+xG8TrEsSzRRLg8yRNR7OODVHboRB+LPGnTW6eD+WIE9LkE2tLp2RWuRfmDUrRN
tBSvEhuCIirR36xKqQ0xl+aHymh41r2fEglcLImXv7Azcge3vSLc5aC7Gtwp3IxZZKfvR5IFuJTL
zqznjx8mpuOzKZ/OmwoMnGsBOzx7H06EuQLELc6czqiV3xF75OrR4qHEcXtayunnLvyU7tN5H6tj
zJ+n5akU/BRKQLUXHuy5djghXeby6H/tg0bD5Ue73Jin5+JruKaQO4mVMqoCPtw46PrcoefSr0h7
QYPOVZivnLz7oe2Mk2vRHMxEaWEVxA01u8vJKMjy4esvs9IZW+YY+/QvvglIGOcyIFADpX+8ViK+
sm+Xv7b8DQF5sf8TWX0LxhHgAABPUEbpwwP6+VtvB8nVRJEgumqTLH0SW0uJhy3/vky27gIJK2Nv
au4AZemEyzXMOcIlpESj8mYUT9ku2LMjJP+w8JZhX48W/VxnP+15sDQi6SM0kQs7Sv57emun+KBi
zN/RtU1/Q3wzj08x0L5YyljSHyQbOgzyoa0gdZrQqvmy024A9nf71j80Zott10W6dlotMD7UIeQW
pxd+3nLPGduCRTgQoStO5vywXIxdC6n3xbt+89hqJVG3V10LX13fkKmK1Y2I/DldDW1r+RE+MQrC
NBzRbmf03Z9SDnSOulN90/8ymsFQ8tRcAOIVYWQY9tb4cHTe9P0ld0qPvlpHFHz15DjioEWqXyH2
VOilUtg5f5vgVV0R7jYDpsYK/fq3VShsZXpEiOcuDeVeyj9R9I+QbE7yvCO4z1oRbx9NMaADA52T
XOKx6H3XcD75zSBrDaMj9Qd/I5ecnETdvOrzUNNPZk96OFz7iouvV1OfJRz1BrY75XuOVW/Qv/HL
QVm3hYIgWvPeXO7dmkPUscRSMCVUMxcIwempen+Ob0+rwP3Pvl2fRtDXNvPLPdDdqsG3oD3gqsxg
RCAFFHOO4UKPQpFzzkHsC9iUheRiMOXvYwiBclJqH+k4FHizW9BQUoh8y9C5iCCeVWyKukUfhAmV
Bh0blpsozpLjdXyfvyfRTKnI3QroNStJZwipwJn0t8Sb3GfQtNx4TkGPvOowxvvx2/nU/E6W9l4j
Typ63jp870D6WtMJ4vhheK+4RKUY84Iqh6m+e1RdK8HYgbYBfe1plsfJDGWC4eeP1jlyLY7zspJY
OgSLdduEDDEd25IXLbgOm/48r0Yyvm7QappIONkcrQBU2dJHqk5sLkOAMIWJCc7iZlxOCzD95g7n
LpX4+Xb9tV+KZFz5NGrzar1nS/3i1HAIMk0FAfmmGaBcKSkhqJM3oIDvwuS16ozv41376DN2KP06
CtgAhCfZVMcfXW8Id3WF9i8qfS3OfZhJCtsQmVm0CcCIF2sp7q1mXg6u+hGeNBqXRafNQBqQU6xc
vdtbcUsB6z62kQ2Ny/VrVRrYnkwa4yGH+B1Zbyp68End3uRHXqGt7Gug2F2dCxC6wZfsjSxAKiwa
lKPGqJ+gfQ2YOzrhGXIbpYTz+QBbkPPsPMii3uUHFzKB26ttwNcAPFyoLdczhYqUCjMAPWRhHM2H
XLEIQEFVWirSUSTBCmn8bKa1O6PGv3J4X4jEkDaLtJ1Yc+Vg+ZQcpsuw0ujB4Nllt5FGD518H2A1
BNkVbHzhEbadEowoLdEGLaOeetRtA/DEFHJbEZei7vEQG2xGJZJFrD86aXTqxwHrlN6Z0MmkXyJg
L750X2z6ulEESET0HPMQTc5DUgeww24g/BLvl72JH/Jd3LCNcu4ngoolM1iVWL6+GcdbwbD6PUZk
1bwWESOJiFg+vl4TkyXhvZZI6WDzWPvhzG85kBNIjcxTnPu4Jm8k73hzpED8nI7BVbyFi7njHPZK
fhm1WnAVffwDiGFrAt3VrghGODATafjwrOtLh1B3rUY758IBOuJSiYh73LeJzqAMVtqYAg6xRoyx
CwoyrSRM4UlfZSLlCNvpHSO/q33rcNepw8dr1h4zbhjjJecOWeB01zNZI0xTb/X0L+SuWbUsoQCB
9g4J4phK5pvsTXTKJa1RMLud18b7tSZ3Y8azXTdUs2glxa0oO5tBdl8NWODpfVY4CpGDH4B3eru4
4KcPo0tHKJZPyhplbCEAW48TDa7SnnSjyKtyutNoXxi5plXJ68UeyDg/q99x0/x/sJknTcwCfl3D
PJvynoUDAIuJ+x4P8aYAcEqovcIgbLOk0MHjMxcRjtQnFxC1kd1a8kzIOQQxuscpijAYUQzQoGpj
qJoiCh7FD/F3XTu2giTmCN+2m5neiPQs8ro8pI5kLK6q0cgXY6OMsH0jM+au4XaZxIbAbHHDJd0m
61g31SGORSkYSKtvwf6cQtmYjNkmgKphSvvrK0wPSpCk+fma494EYUeYdheSzV5anNm0YvQ9qGP0
UGeUaUckbWVDWdQgocZec8JH4DJ/80cFYc2TUjUWja0Z//2XBdaWxsFOWske8qqmQRjrLerMEnMm
sig+JDG1DXMnF4wvNdEJLOem4Oiy85cgtVDVD22SPnHJ2VEz32o5ZjWbX0CoB7R6Ykx6V4vcc9JO
/JoCR3H4JNp5SmJrGPe7GgCM5LYTIAb4Eq3L31lQxHT7E77cuebpT55tDH2haDmdkkHWfQvAH2Fo
FkXjlgFo57Frow7iWSE9W3DumQozSjuZJM8j3q0TErNWMrh3eSOut5KTgrmDqtCv7N6TQcal/oYe
1/ZH64P9RjWcopP6un4KkOIFxVdb6iLXU8HN7K1/BxIZ/nn8Gxbv1+N2b3LeQrQ+7XG1MM98TpZl
nqBNR59fN8Qupzl8t4mg5yY2VMromjnDOUsj1QvwMwb8xoUTRBwYVq2u8Z/ZkhQeHRGjcQSS/6e7
992uKS1VhATCJlPhso5ptZoU/r2qpsiSqmejQtunuDgDYyGRXGhyYUrXl7oOPkVBprJ/eT08GMjc
lRegF84NMeuwET7E3neCUdbCdVLMczlUXDLwASJzDpWNZuMUX5SYfZAeEXJ+p1/FnuigfaF0I0zh
jmbYbDNJEQ3mwZo7ZMSRp644x9YS/wdaRfQLTUF5EQdfMgX4vjvvOK5bKlnggOE7asL++rTdZ+dg
d62tHfK7+yCM8RBGFgI6nPn1bpnrzZmkFAvy9H2QSJHawMHTAG5hLrJKMskA8uiHNad/hWF02mpm
3Ger/Rvyv6z9CSBzeNTPV0lTG4gFfezm0Wea4bb6Q72UxEGYPscc9mIPBWVNKOP9BrgnXp5sxOQg
Uu8IVp38gzeowhmUV4EF8fuBc47sYH/uEv4IgfSNQN28uE66CHwliP7OjcKePWMnuyNeNnTK/j51
0nMhQhRTU0dkD6GCfBKb0z3u9bWEVy2U/nSPpLPt1Pq4IBSVfDWvfrzIjydnkzriRV05YdqYZSx9
aTaeG4YhojO3RsLc2KHKo4hWv1Wr+MURqvRlC/uJKLv1N7mEVDB1yL9V4iJAg333qkCMEBo7bVlB
ZUMI1r5ulody+X7D40Ac663jrGAZSdKLWWk7s0xX3agg1iP5/LH2ceXtfY4ynzGvulSjaMhkXMOu
K0rAbY2p7PYS0afQBzhg+bInpljwly3ZKkOb4oDrVDWuSJRpHcaO1/z2OPgolwOVvjxKXT0VTMkc
FFbTX1Cb9ntdC32SjWkqmTNruDSLK1YPV+ueXRsIC5AkRbA8rk6Q4lnlrI0fBJd//6J9dNfKZQ+Q
cno1WUFDf6EaLSE+aPV66zusBMJkgzq8QhZ/IXdTvQdduwprYqNzjRkHZIhOlcLHbnZ54ZMCiP8s
Fh5GHjDUcRTLea+3bpxrG4rgMMPsxYgCtWt7KPKvG8cg/dg+0hAhFjyL7tpBAcfGgCQEQBhAZUVg
7jLpoayTi65C1KUB7jFr+C27QIc4O550+IC2nnrjyyRh1pPknvEUPNuDiL1e/Zbvewt5+u3lM8Yw
jekQKGnkLxGtmSPL/yqU2y1L1EnDxq+NUOS8cId67I8wdQ57jaGnbo7YXcKr3NSAyDu18O/NIPWg
JvziGJssMI2sPEOq8T7xdsxtIvoNwS3PjhXG//Hj9RZAZUTmPfgPT/J5XT5yc0N6zjXSnxxZ7Rmi
90GNVjRDUUbESMqZDANM8C5eOnk/TSBun/S6dZF1KH7khaKyKVG4PIVNGcNAnRg5J8aJEkJVtPuN
NtpDfzDCnC4O9MVHlWkl6yCunm3Z2QxFVD7Qu7bsfp8xPwufF1OQIyUEyV9GGG3cC01jGtRSUqOn
U0BLvhL0VD2vpfkHO0D5/RNbX/XtKkq1vvGNgcuv/NOF4KLImd8va1IuZkDIQOJZmTVFyV0uMtfz
6MWY+L58t2sdrbtywDyrr3ucgUAYIEAuulh4sHkY+SyLggEHIR45ojv/IRSmOYsSdxhb+W3rqTV/
ICXTYhDRYTPj6cy5CHF2Ypkg9H7P3TMH+JXzvY4Ms+XSqtfXa5O7EUPW+hz203XkkLMi0Bx9gYlL
+WPimIb1hX6G29UJfTdNcIeKcOCxG0gECZyF8w5WJUO86GVb0hmjxAEN3MH/IpxH6HRtrTSfjFj4
Zw/ix0xDEk2J8pj9fvuMBPXL/J6K0aGKUxR1U5BrVkVhS7ftZqdLac4aYkWZZYi2O6lUXyM4r60a
j0gT71QNZsHLJd7Kbe18fpJilImxTQwBU351jvn9+FKQiFXUkE4TPWtuxhy3/of+r9xp53Qj4XfA
+QYEGx3tkWyGeFR9vE8/8Q5qaguzWVro6BsGTETQlmLNRmnhnn1RY2UEBqpoS1ZafY1WHnieBE2u
m/NLgUrhBoX4jQ5UaEW7T9ZhPw9lX2lZOlDAf2TESgnMbvOMkyLr//Fl+v30Esmw+0nlAMFbI2n4
NSE887A1D1kzmKRFfHlLeTcFbpOz0eGRL33gX8f0WINYOUKugXTfLpCItCIJM5zX/hEkk9R5HTxS
vIwWqW0eNmrXBM+OQrYhxZuV/USgEZKB7GB72UmhyreObI4OfnT0dwaEqSF+N/QlW2XTFQRom4E3
bsyiRbui3l0QtkjZPS9GCmTLJySkany+AjVl5+5nUiL95h0cE1cc/49gAXN87zcYzdrAzbX3CjH8
QqaekBwk5uj1/m8m1Vbas3JLo0WLqfJEYDXNwvSF2zJdpY5CdWFc00OPcxhlJaWqXMBnP+yBC3a7
PjKBXGO1G2h3pCVPElUxlTdQt38/XmY8MKgILCE0i5h+38LNTSQ6ikW04/7DOr6wn6Q8/ifPpEPL
cZPLPWtmN3smdPyx5Uo1+Peq+glnl9BJYHOvDOjeMUQLdP1jQUIzxT2RpV58OCGExELv9NJu1PuL
Q91ZTVmjI3DtxJOQVw7stoJEVCpfFzWaFbDjm32RnhPUojxD1eG12kExfiU70OmkqpULkJSGHuZf
IC881DQFX5WA88cah13oCUo2KxbrKf//32FkYFqnpWTciIZSe2U7yRQHRp77J6shIxv22rWhf84N
Vq2kktKyjK0etjmnNRhCrDKorFVk6q6SXyOsUeSGeFJ0dGzp3JW9S215IGI4+F0wghBqXGM/2ECa
eEB2rHgRzHRiHZefGqI7mcwqmmDxnTMN80zyIlPyWhJvgxveFE32GaRL6jp9LEKHkwiVPnbz5K3L
d/HsYgNfR3a30FQrxDAAGMCEzH6t4rsUn2+JnGVDT0VBTDbXZGE8W1COIFEb0LkQ+d150FtCg7mx
V9w4ZE0R1fv+UNk6znx2FJGks05YMuw6YMt7jtdxXGj5msI3489VEbPzYv/sOcb7RxsSfqcd09Vd
VVh4i4jssqm7MszhqwUCXzV21Y9Ba7+F9V7s7t7NliXCBFdduLCmBxBAz4RG4P73yoL3vZTGfiMt
a1Ak5kZzuDz5T6H9cLPqhtZrjS1015MyYDnHFGYs6dlQaBKUP2JX3/rpCZ6SFeHQidgS2y32VABm
3GN+klsDJlO9uFsJlrrIXOWIOEmZ4gJW46D+Tt5fvOHNQNaFrmIwM7exbH8HFsJ4YSxSL+XaBOAr
rah+J7abEmwMfhWYi6qArWObiFUp2UjFPIfJJae4ALCh+aOUT0M/nHeCZJ0Wh2gwVT9uKVFMlrx7
Fji+I2vxtuiEW8wTrFuLenZrKY0wOaOnd+2bWW27w9IsxQ1HiJSecs5LMW7+jPPSXyv6QSCzJMFU
5FbzaXl/vAt+kX3dpz2GbXnhS2WCGTeXkl/7trtszTJqIC7F9Rfkv3KYngoXUYrOmp3yUpKxgdVt
4b38gkjfPC3vBcvtTWwkCoJZBdAU2SuxE+PEEMAQHFylEmA8ds3UW5F0S2yPqPjdaF2yLN0DZVzf
ClYA/oaqdnakxoNdMBYQurhAFGHMuFukHUZ9w+/hpTABx0et+sy0W9rCT+VBSWG+n7NP06i2tz+O
ogDbrsh79K9ri4I9GFbCT55a3Aj1wQD+FA8Lyw6ZOrXQsLdNFiOiQgESxif8uTZlkMh46jE1Usm1
TPEeN8XKBpwZOvMq1S6pvjoQifHEABRZ7joA4Ek4aQ3vXTgPc20T5tuJJmewxdMKKYleeXPnhcGf
TmLJhVLQ89IygF8PxgwnCRkABsYqhliy5UOzK+4kTwMCs+hcPzLsmr5grzll0Cau0n8Xdck/LqPI
Mbos09Q2bcyMRCR7Vbj+zKzbFcERxf1Sh4Myr38vFx0ZIrXdq4SDDYLk724VPx4UGI0MLv7G6E1J
jzApt0o6UC/OPYe67fYPRTzJQ3JTzN4j8khNvMBp5KiWtPdxRm4ACXYyyU4AqCLiQ/NN512s8Ega
mD7OfYmhAZc+7ixhG4xKkkePKIYGWptJ33IhNYA1HHDF4gTLE+Fkh+ACAMeKCOFGlxYOZixdvXzA
NJ3xWNg9ehwOPZy5BbtgKZeypi46GPjZOPpNGusZ02OzlKVzD3YK0YV9wKeERwtZJaHoSAWIWEpD
Od62MOWM6K9bh4rn35cAbj2Gf1Glh1YwoQwMmD/CyUE2BYJG3i4XJyQwo9q1O+t4YUy9ZIhUjq+t
opo6Tnd1p4okzZo8PpCHuAuTu2yb/fifs5YDROYkvtFRV67Y/1EGA+3d9A++ZWG1SQT7KuV78PoO
LprhWI5HoN1uEkHN9dDT4PsVv3x9N6QrswLI5UTwZoGc4VVjdguP580To2fHu0a4HiE7IgV5SPBu
vyrE2nEqcRzi1TJzwDYZy/9RR0lwFpq+xArejgHGaFNsNPsiThX0aqQHVo+NlN0dsCR/PCMpFySv
aYntuCx4KNIpOERwThUHnC51uQZmjBpv4gPXaPxiX2eokDHwG7UTCywktTjvTraPe/sNbW/eQMIn
rec45bZsIrtNxz6rp1f+pZi0AaY6GEAY3NnsTcO/cUTd32ujlLvdzW/3F7eIXnNLmZevugRgKIcO
H/bPBHI1uRTcE6AjfElio1snSRh719mpvvZNuerRrx2ZXF5/Pcl2D4xIrD4FX2F8aM1Xf+i7Nuqd
fnv7mnIq71e0dbJutE4W/KbkTnjNGf3HAGySERTki/qHuvHYEXCclx7PCK042hq4FGYK0dUNuJUB
57356fbXshfWFWp98qQ5Z//nOCEbB7E1WUzFEMTVg0hd8K/U8Exj9ivhFbwCzCxRWWROJjQlO1OG
tTL+x8IsL37UsV9Tp9Q5yjqJ13BtcnFUPnWlOoasXQebtRIYaP127eY54HU1oCL/kxnnGEzii1Qs
V7dpzHSIcqyHsyChjwZ5Mg24fUTvK3pQkSaJcKqP/WYbPZoQ8baeB2h3I8JPKnCToirAYRzq5do/
Z3VkIA0PJPPjMvfgVoegliG/u6jW3G/SCAZmv59oyh23QhMGAz9e/XyUfdD+iJK7gdWlF60M4DFR
/S/IiAQevZvD1RefQcylhatnIcj2oo2ZNwF7PYh0yhRDjEli3CFEY+xNM62E13vHbTcSsH6CvUL0
4YoqAlw8PAGGh6UC4q3VvHJdohmsdzREldIFTgDGczzjowk4g1uQyzY18aGblUDb2VtlhmOj0iMr
1Ttd9AQHjRfjsDPjD6e4/1WuxPQb7MOMa3Hf+S9dDhPV0xtsx4xw/rUmrqp0j+8TlxsHWEhjzjPA
RfSRgnm4iFuQL37QbHd99gcpaVRR81GKqSHP/Aafr8cHVmfwOWd58xsIvXpT6VZ5gi2Pv1V3xNnG
u4tl5m0OssF4jg8PRB6AgyAN+tmxUeK482nQ7Sz9vxxipzXxoeoXxWGFqStY59rNl/E8p4kPZ2LN
RVR/+6GxR62UvHgWXYMkWQw5QCKbTTP21kBvHbGFP8X2ZtTc44fousOGMphiYZBIBjMNJdxzWDXT
re8+XLV7cNBrITDzrnjAGyRFr8HRL4eHdpXopxlmeFzj+nQSNJk9SRuTudCNSSbHsNzRtq8hS4Qh
IZ9ibIvzZBOkyPax+mrskBNxnZDIWA6nI6DQZAThxHIg60KkzOd4vQRRtoawX+1oWEW35qA8szBf
RQ2hVGl3jTgraML6VVrXdejfEkVqUx/fbUV0FzgP6Hyx0yKtpzz7idKKGNChjvn02TRUDxCKRIpq
IPmZSPI709ZAHLRx1UZ8+GfEXP0p8OuBhehUX76JLgN+toeWHtnez7fiviya4TlkamevmraAxAot
tf6U4XSIJ8ntjztxXrQDVR4hS3lAqw+kZWQjdycWNEWIoCeOJLagFbjdboNGosuvGXdDKiTNESro
iQWrYXMtpbKVbLEiEtPswCp2krpl3CD5cqWb3lzR3TPn8LEaG7EOR3IEw89yptG4MdJGHf5++iOO
dWz0cwVd1U2AnzGepEi5Td5ub/k4T6xHmU6z9/sCXnh6HSKYLwyt1Tabtg6/XWeH5+rb16y0Rrwe
Mz4gnJXkrjyURFyRvlz03+8E3d9A60JSx7wU8/393KKqCchKiNtM1qfEb6nhksIzpEWHImjk+VSN
czJUWn9ScFpd0ZwrmUsi1rZjgpPl9F8xRr1EsPajc5bG3RkOcleNJu9F0YPDHGi7FYv3qp7hqBlO
ghZxjughSuET3+xjWoi15NmqWkFcAcfOc13U8oZetB927sWQ61r0/pWaECDHYzzewSJADpjsEE67
vwmoQ6JxHlRycKqjsePjoFVEfjrRPnG5aBQMgKaSjOOwp+OiITQScFlZfFbET1xS6C+Zn5z6IoMa
RffXb1KQRvoZFaWWk3Jmq8Ps2tVjjdslk1KoYt3Yiu3jFI2+mc39l/jYlkPhHzB62/MSpdP8DCu1
2XLt5VduULy/3TWCwD5maXyANdu5EvYrdbP12gklU8WuG1WyhPdtbUSLtTchFbAI0NOulwPNlbK1
SktYwcuvNS+tyGQ7ocINAAuMesTvkrfcWM9PXDQYnpmuS+Qxuedx5dYE6kh+hdOg+BAXupG2td0F
ajpD76yARV5zGcW2Z1otcbeiXl9BbaQy2a1MAQQDMuXO889+MqUPKNlPMtg3+GhhlDB5VtOZH8lE
xQJTfs79zc98kUSTj4l7O8aYd1RiZAHNiF9D6zoKKtFsai2AXjsAkbP31+29suqugZOUM/n3QEdP
COoSWZQjDO3wYJETpo3IBl8S+bcZ+1AODRSAYbQL2klrlN6a9xJeVv20peyzL4nWBJGrEzbYdxsH
Kwqwtr27S4fc/mNPU7OvN7GLLxWxl/Gr4IaYamhGPE1LdmsBn8ThPdiB3ec1xPXqOI2uc0zQ/qCj
4OSJShT9nTH5eAAYTkZAwI8ZLgdMQJcsPbuEel8SSYYuj1Jz8amlZutmphtob/JxPJ8oTFwt9L8c
xUxHw/Rzi+KhDhL4CbxheMNxABRo6NP1wyU+c/8R+aOcCj5XL0GOl2lcXEqZjXKMyvBpoIBvLjRt
UEtoJoLhoTtsfbX+tCT8bvbvcFdPQBMZ/VK78oqTtR09H2gAKhOJrwjCJhMo8QaOLQrc/BB/hUQI
77VFlG+6e6nvl/QdmjGIJUFfvxKHr5WJUT8aAD9WNrD5jG3nCCwWYTmWK1O4Gu2IHfrLCvJKUd9T
ce0AlTMF10jDFIsNGfi+dQPgESAFgaxKN9KDswWIRbmyZGAcI0uxkAXjKXSrEwWZu49HOFmSrhAr
o/YEwNekM255lubg0TyXrCeqaOL9zXb8VwL1BQFip4i3+MSvw57/4ZYTnIRuaIRnqtD+31HM1oMb
cNBgaBprr2AIsIueFPnAV34UFIlGquS5iwY/yL3VNNG383MWc40SeD8INKfN29aP0fQGh7swC8Gn
FH2yOFAZuyPklhSabKVdu5m4PSb53H46kMx4plN3010P7szArEQ7ToxhgCB/gu2+fFi495TLVpJQ
dCzbrK9LhnEfj1E9tgOVo3Ls1VjOZLFwzr01ikfR24EOd1hlqL8LtP8WvTaNVZ+JL8yGNFPRWsBv
tJpx/H+7QgmJX9vwqpoQZ1HjT2pMidUNJGgABbHk58NH0WYPuMdoAy9ITWxCTa6omZXx9JULi6nY
vTEW7M7GDPjWWIcD4HUP0t7AgD54QfYTf9vyxuv2sEin6AzLTXMlv+02XZgmOHSP7haiNNefuKtP
Qr43Wh38JusjlfSmNkGS4mdGaoSmNti5uUbjxS6PbDilGPSg
`pragma protect end_protected
