// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:54 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
WeNBnEBdl/rEBMR6FhIYqj5z8aTJE47BBMVBzs5bPw4y3biUGPBxqTBL3pQyySRh
uJsNy2XGYaZjV1Q7uZGjgT7oE9q4ZGysCKj9hucNrMhB7tO775AvZ7ENc1NIgfPI
qqIs9Q2kBSPzCxEj5KWOZyWL3oBEEF2ehjWbdMSC5Rs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5568)
1SQi+jFCnc1ofOZMBl078NgJI4o08a0ylFDiFYl/L2WCF5IpBnJ0Jwsh56Ynjde0
agfLJJ2/8mHwduF7dk2FfbSrUjQ7iE1I/twxOwuXkQRM24TVQN7BVt/kA0iQXhEM
6tjKEnarkarioKY3jpKten9L6FEJmQSq8a0VKF4LncU2JC6tgbBmZK/wqwzRV8BI
4gnYH4vMd2wX/39dQu1yYUTh56meFjzjgLMELqTDZl8LHCT/KFOauMBAbysBBZpp
vaRBKYInnUsjp4ZE3LWVp7N6oZ0/66D+Uho82W9bTX/WixDDvQxJtvXbPYkm4DVH
ZRjtdEH5+OV5yTeyv9qEJxoWBAz4bKJS5fXJHLWlDRlWKhsTY6mHOcwcoz5zYunA
uGCjWZNqDRJqlPAMtA+UsXqHk3IRqM0WxDMrxGRKjD7c+sznkWe1SMafslWnH4mN
2AiZ1El2vlOsUGRCAZOz+1r3CRenNi6Jrh87b+uL3WeQjivvltWoI9cpOrOJG8WM
H9yuCcnWdP+9ErvsMFhp1xU+vETjPzoDypEStg8cK6SDIBkRqGxbZWsfozYbQX4s
iGSIlpHffCzf8L0okxDAh0wiMDhbktXk0D2cTQJbm6pX9phdBAXPzbXHutywH3TD
w9xvD+lcnbbgSo3mpXgW+s8VNXI1hZd/qc+buKcSVk0EC7dy6nO9gSO28WKKEH8K
KiJbpuaabPmQ4w6tulQDj4XQuMZjchtYFRh0e0vBVyOSKlmop8PqpPAx3v1HD5ww
o280qtabOcu9MSZ9sZwNtvHINkiV/WL+2nuJ0zX/t0h02qkNnuAYM8vOqjDSPadv
SXY68Ukq9+M+B7KhpU8pcbzLYtRcxrBTDrn97Exfl+BWNx2nVn/3IaT2pZS2Ck+g
Gn7+AIBpgTkua07WD/6wr7OTUHz0RyxebO69X32UpqNjR3Fe559AoNYlK17jx94c
9l7Y0DBieIoTvzvPiFrrjtBtQWP7fHtSAf2+F1bPIgnIamwqVDBQQLwO4UK7+ap5
+cZmQtNntUJkDzsEpaDXJyygTYydN+wyyym3IKpxKh/po3KoIZ2MlgmDJ5Tco7Ok
lSV2GgMx4GvOFGE+UMNnNOk4dwQZM3yQ/IBLnPGsVwoeez40XIvh+X5vZonMCPGX
yfC5qPaav5k8WSs5FhNOLKLBxiO2seLc9+BcuFL4o2AxVJ12FcciV5F/5WGhchj+
zVt59pHBCSx3c4KtVJ2qJCdvQwtnQg8e1GjQI+aWfxdZWu82pHhW96ThAu/UPTc4
IUHQR/xUwtCHUitzJAmCeotBjKoZbb+Genngmh1psj+ePLiLDb2I2xErFfcUsIbs
nvhPAWRcsP/gs3ceVySJvUQDgRj4l6iEbtjPRx800HlTkvCCLlYHwGA8heEZRsSu
WT1AGG7qybAP4cUvqnZAzH1cbEH4/MrNLBnhxDFzQn4efxGFKx6+38roK43nhE5s
P5syUkHCrw1MwlmTm0K81+f/mCcIu3C7UgFMMEVUuZ1SFfpZxTdMULW8S167gLZ8
xCLRP6PWRpl8ZPR8Q0ftuJoJMwgPm+fNiE6knlhGwHEyPxNysFTTOY7xKuehldHz
5kifnDyiJRG66QHnGLUFgcmJSktQlIDaZhRRkFGnN4QYg7f6Dl2LOo/wTp7FMM3g
XV1PghIerKG2NKcpGiX5kZJOS8TwqQxn6vVwR/LIQuVJrM1mAPUL73LXfR7yXDoD
w4lzJxEy4h+4zYpSHdRy2JvvgjhDxTK9cdLQsvEpE6doP+kNtSnFNLYnne9Xn9o4
5ylkfHBljXFkJivIviTLViNSUfmep3IPvZDMLGLOLSi0QJbsBNa6wjxXlabNrhWa
CWXjFXGPJZL6/dcvmnhWTkURYlqGyj5O7qHGm6m9SunEiHzS3KQ5gfj4Io6s1iA2
e/qqMLSQQCH19TqK2U98b+Mn3z+NulZEBPgsyuyB5HABHLGigwTmyifOOGMaF+Zg
BcVEfaZyeaT4gDigsy+5vWHZm7icK8YITsCbbRTSU9FkS7hmSwfrzJkPELZayPrp
EyhCkefeNNm2/pvFS4RThJWmwezZo1BL1CTTGU162Oxfwu6y57ERit7q4Ssd003h
1G20wJ4q9pLiLVYmynX7KgfXiyzjFt3XTCDbosbwSjcSMYiIqz96isL4Goe94uIs
Wt+GvVUvUua2a1/iEyhoIlO0G7exo8BJEyH2zToRjXRL5W52EGIhtZo3AjJ3PBSG
r2sd1oJHI/oEj7kD8EtLAyhJcEU7omR7nP1zri+kBuw797KLRSw/sn1YH1Brp/t6
GwJfyyRL8BMZAHj8K16u3C/MgvwZ5tgs1dXWqZyuL4W+HYSqMb1I9XtMaqbXQi3e
1SgyDVZqq3ftV98Qa6EtpZIvGzaV59xa4bIBuFF0GnveGI1yGDqXR6lp8i+c6d5N
IYJtLepZOIWyxbNIDckoFBz4K2m3RFQKUH3PhIq9MlTO4dCVCnt9jNPfFnXSZRoo
uHrsJ16ONLZLz/KZVf8+CD7RsXwiheU17qcGlfvd6smwJuxg+58qTjTDHvooTluS
iZW3gUOuRYMUn7LduGSFYJIxmR3FNv5Hoodw6NCKyvzsRSlXCZf87IdRiwe8t+Av
hRwqcbxh/yv+r9tE7m2hm+ZOnS787rK3pyjHPS6rDF4kcnV5DqEQGMNF84lQhgUP
r25oRdbqinZksLy5F4qdqa+OG/vL92ePVArGmPnlm0NQZZgUDB+vkFpzElnzQWjz
hfIP0miA9MJnVdrmCiQX+iag//QuV9spGex9LiCyyld4eJxFYnETTVgDxHxGPAIk
dCXY7AcmXtJpipihSp5lz5GAPC3klmdlUyJGrJnGMT+L40PSt+05sOvmORu9ZIDI
ZtgUAELRw9Fha9IZbSCESZfDBm7YCM7FtO7VNFmcQMbFtfTihH72IwDrQpTxrjs4
fekIO7vHho4Fv4BF7Ut5yrpFWJMMD+gKf/HrdjPsspeePNxXMwQtuqRbOkR5tnmC
hCx02W4GrGFmD3HHEmk+GQyR7Eiw+8UVU9xJlSBLOy9d/zU7Jrau5PzMly1ae75g
Xvn02VbWRWmVU+P9SKfb57ddZdedsrBq3GszTOYAo2x6POlWg3NTOUga4LJKA2sx
QqvBTYbZtpyMALWiP9YK2ftqk1KG8R11aH6fFFCD0MZ09OedarB+IuEZSrki5PiO
8JORg1JTArYwNP8JnrIWhaPz/3RGWp+SrMInv7+IeTf/tjOYxt+JMKCDx/34K7Tp
QYoz1Rxk4ZSWBKX6BcU23JXaJp2FJBSgIacIXDpm9j+TM4ZQgPGagkOqrsW3F/zS
o384E6w0skpspOgMc1gJfbl+QxyJHfhnRHRlH0qUndJfgYPpWk+HJJHdRnVO/oIU
0VnoNgiV45KM+w09ZaJiESCPAhfY3x4NEhddnTdzs3BPPKdAdyTj9ZdT1vWgUBEt
a5pNV2XJlop2iPUfbHRRYU1teYXt/kw4uQnX+Ucv2ioM9grxY4qTGD4Cfsw8sotx
XGdbniK0tY8K6fDi52fJXg4ogpGS3y9wwEv+1qk09sqt/hNdi/8L86MwqPbbT2z2
DQX+OXNoeY6UiBOTTKONYj0TIV7HXFKSViekJjw2H0VDp3rQ4C1qfX9j/avEj6Lt
WqzsUEboM5j+Zp435TYgn919HZYuuDSE+HlATW/79xKPoaUpuetCCYqeyfZf2y+I
M0DFcBYY2l1p9CHcVXPHMqyFkwp9XuL5m2IuxzkiwMuKf1DeMdlGwT/d5+ORuaps
5vOyHxBjp3sngFy1TU1nPFzypNJhKSaoQUSs3w4tysoVYZrAsqi7EctumGdBiIlO
GtfQHnGdI/Iax2cEa/NomsdcqltjHOPBletgQAApYYVn4Tg1CjLHGSKqljZd+UMA
zYX2kvudhZRBrDpCWpogS9woXv8Bnrc5F9JWUQYbbc7U2khM2qzp1LB5QgDYvfhY
WTvzNULO6+dpmqtLtngl4Zioy9dvMxDmHDp4XMe0DB/palvI8vXuH6rMAI0AamYM
DTwJLrd2KCQzXQf3BpTjfJw3t12je3hqxjR4tv+3Auq8fdjxOiNHa/6whSBfBuox
9bGnp/ijcUHTrtfWc6nmOEaUyspKG0KBNSyybDS9Q7SZT6SYrCTZ6i1al+iBhZKC
kZDbLThgK17u9zQz7y5kdRLF7+3388VJB6w4qpNbfMzGwgopChNIcxm8O7quk1im
74G0i+KpdFoYUXwBCzhSIN15amiiS+2XvNUyPlt58XqhdSsQrp+6V826nclWHtYq
15v6wub5khJhMQg0R5axbjl/qXuKnbJ6b3cFVuUdbK++ccwUDy79wHTCaiIsYsVa
US8GgBvRcAixcwK8b2u7AjxmmOh7TBTi9+VQVupKeUzQAz+ANLmAUXI8j8sRfxRf
mEbvxUO3Zr1OKgwL2SXYslDIZsyZq1eOZktfTvsEWg19vrW6wOQMjnpjmB3vPstj
J1zbChawzSPz70qoLidTR8iNQ6BTqPvkAO+WmUxw/pypz5uiuX+xFHLZq2v31Kke
kls2i4LokDKxu3/D7YxRrolY56/m4SqleDXN6HEVTUuWj1E4GmaxWD+cmDp411np
+ogscO9NrB84Y8IyA+xPRKgRJampll9JuqAAbIzx0sthfOGNtpyoubdmWIMQ7u8o
cC0gt1LNI8tmkmq2UvTgnHCAhSoE4RRHP7Qqz7PBdvj2ypX7wnglSS5rccTkpGh7
jV0tw7KcrmMVNcwCUpZlQEa47pLT0ojYGNuAy+C7hktKSTQFfwvCYKZ1ehbm7SPO
GoToSbyME1R2mFMKxP9l24SW5CbH050AeUdlukUNcuwQ5NV7YzVJqWDnYW2P4HT/
Yxb1CDO7QCCELpyundG2NiMLNUSngj8qtCtJogpKlGOCH21hkfmWSyfvfwfQRApH
I5KAxYNcbvKJ7GlNL7b8mkrWonp4teFXc5+9nyN36nxZcuRUQ2F01kYgWlEI349D
DYlafurH4VoHruroShHcQWpe0/R1mBXXU51h3KL1rnSUQna2RU5xVKL7ouoE5+bP
BYEgOMEbl4yGD8uYIsCMrPABfDqpkIdoqCPxyzkCf6U4oS2ajiyXlsB8OUdpzFXj
eka6aaCKGnIJyebfd9vSpP4kYT/Ns3YB/hOqA4J6a5yNp/WIpuJ4NHbfbwM7x79T
bKE9FWVZ9ZjVouexbhYJNUG7kgJvb8qzyrmiKnmc4P5Jz5eMyWfVa+mMOCdxDlXy
yofrKuvY5Cc6QXPXhYX4SW/ujKHzKlLNzptxZmOKUohWJup8Jvf9HyR12QHE7Twd
fqwQ3D4pL19bFkmYJSKX3vFrO00TL3/BKEDXqF4r2jeWyD4fgUvSPHPlvfN35wO5
MCYrn3XT6DpuJ8WU2+9RxQWk8pWoocTy1CltwiTBHtIGsanKtT+kl5WoRfyNZ+GG
wmLGbkpYGk3OO4loVZzjrbW814CxOFNHjhzPPTaJPNgGcldY02DvwNwt9nHM/sEI
Wa4INFLclReIMJN2KrT0acqNExQPADEUgu8cfjRtC3MM4v0QvRWsggdaqRolNw10
lZuFfrRa67+SObL0m/nJqKKknNDRsRMqpb2N4LRINJWGbw3ImJO3I4udzw1T2J7g
A33Tx8ie53+fnp9lAqyIGkJcTsOcEERDrOHpImtNPlWReLKGdbXX97AORozhxxpf
j7v4yovGp7nHZ09Oh69sRSfCy7F2lMq8nSB9W+vFT4wfR5vzDmUof8TcjixWDik7
s4jOgdtYhzI9F6bZJyFnHit8kOXnxvMzLs6q6lv3BUmlE76Bx0TvzM8DqvPDOiym
GhPJyGuyYZTihGQBYXkv9jfFFEm5fcKVoHos+gb6S26xotFbwID0VfOJsDb/tfi3
dTFyx1lGSVU+70vJ2PGe9vIFRgBJSU3gwj4i+3dpq5CLDBQzdteu8C6i9UNRyLV6
b3w4HPQhKgKZ3WoIQBcGZJH22qDoqKs8X+aF0A99fham4ctBIsboGuLvRPf5FV1j
daAj6fQfxa8CqcDSbvtH0N+zzS/o32m2yeKN8BWqs4pT2x3WAYOJahZ0KjkY3j4p
uOkLJxju9R6/OPMAhgpf+4e8McBMa9zEmQQEI+G0z9j7Aoe+WUjllE15cZ/50+YE
uouBx6e+Hgn/ca0bYX5O9hVyu4DiwShptfDJ5lKOJO0XlSS7WBlm1AKJ/YDuHEdJ
ULQELnEqi0FPJBqYeYDYUEWw0s302Y56lMcYIaOQCj3HcMZGRcgm/Xcx5aPo9q9n
4nMqPsIpozbi/91QO4LofOjUv9ZvbGFePAhkDy/TV9DKg/Kh445sToWynvGCW1LO
se5G+cnIbATGU8dccNED4yFOKh9o8IDZg45vKGGDdUAbg6MPE8G5zenxbuB1EHiW
+7+llS2pYT9Rlgk4qJIhfQN/0ImcNlS8ZYv8KbXjWlwhb+mGRGuyMP37oA0s6sIS
ysB0uQLgEcbPVLPZ2cTf4RjCm7y2r1nC6XEB0QTZj0Jos6X2NUBt+S0bTzgQ/WAK
RvBNBeKJ0uT9h49coHhv8MonL3TXyAVqiDAoDFEMm/kB+vWHInrA7LuPgchu8ZkI
WUAoXi7dp1/FI8bZQQyiK33N4oy1j+kiZGLcJIrFe98htmdLcHMmTuQg4bZe+tSr
cHvLh57PESZG0AtgqG6tfo3cHW+2XOX+lyemH7Ymcq2zb+XFOOPNVZeMUe0WHMya
u/++s7Ru9wLNf9PNlcE9iw4oDoVEe6gHg2Yz09XT2N7LKFE//p387tnjq8wK8yk5
kWlKBN50jXTaBpe58FQCDTi/lh0XZKx4vLzElObe0RsneGcr/caLT2bp1TSdqeG4
FTF4CvAbZwZnqWUXLEA1sKqq/PG76Fe+RscWFID/A8PDQQ0IBcNJwLhiifVpIhby
LcrJHprFQ+voaxPvoKNKVqk4GtOqSqRRklpBOZ7fro2FaqpOeWwkt9MXTWCrKl2j
wfI7PH78ydEv2NN1eefOsejW7SOz/FmQte5hrZNJ01/pG/0Y2ji41N1PKtfnlFLX
ZdOL/pz0yFLECIG3j4sztN85ifeG1ZwIFvg00L8ZsiLW7fOkhePZNOProvW8MNXA
wTyZKtD9RiN9C/Qz3M6h4CRtiAfvVB1lsPG8kaxYrYNdwIok2W+NjCBDG82FrBty
7axWCHgKbuABxBJxyrU3+ATW5iTI52S24W2rKbqMFwBNGyxzwF9EFVU0q5ptwH+E
265vq+RAE26m5rylncZKM5vhxU20ERQRUtYCW7oCnoS2mN5dUfMmtBd3/GDJfNEI
E7fel2EjjVV1CdbO6llrXlauVY8yRpEiSULtlniZ1Qr/PwiEN5U0ImK3YZUxq9dV
XUiYgGCZOKREaertxlqKvJF27ONjcmOiMwVmmv/ANiSPdRpQ3x5VFp83bnBCPQHL
`pragma protect end_protected
