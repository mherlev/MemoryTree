// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:54 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
TzksbK/EJVxGRQjiAqOZew94gMwFYjmMJvykjm+UA26KXHINFcdIMnJ+VkzBEceb
UFKqeAO9K+ZDjjXyQjBfc0WsQzKQbRNm+aeGCAYkU4Ih+t4aY9ulzizz+shrlCCN
g8vMqFrCCg1iOBrkMmKeTqP1Tig1lzZOS4M+tpQvT4s=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 18896)
9dIuVj3RvyeTJdIFRFXjEC2lS+23pn0JB39ru3XNDp4eHhW3xIWKUYyUEW9dBIO8
EJPsKXe4+H4NBLF6g4SBY+uHzRcY1DHb9spTEHNV8jUNTTDAmdoPVQPUNi+FPdzW
rETU4MFJPBH7qDWGxiNRKe+Ad81VffBzmDEETasvD4UxzV6SDUBYPMxkFLJ9ODo8
QfvcLQ0FBQfQR6A0OlkBRMggZYWpgktghz4Me/iLTlL1dbakTJFJtj2ILNcWwEum
+a5aTuTTIgR37rQbADHzkgQtI6zni8ZDntIOEAIg13n4s93euxL8eUkFDNmXJZ+S
0if4IlvG5EclZtsSVsN13OdhEru76W01X/gS/mBkbn/3ohDxzSHeJOkmIPNlcvcx
ushTl95RNyGqKOG8VmxGE1wZmJkSX0BQxgqZ8KxUdaVBKceDiw4UyL9INEMGEfyh
vLo8fHL82AeiW4+Qk0f7tMBH5sZPofCJTzYBugKE9ukjCFm6Okw2VDy6uwTDNaJR
N+ZzNLSYEF3aPModv7621p+QkseozbxDCv9znZNlrA6ftoSLJ/v4hIgVnQq7H3MB
3Z6uwPCv+9oQhjIyaFeu6JHzIOlUbGez9RrbOmlJPVwdaXhw0U7XIgu5sP/0VGb1
nfag217fz+vKqAcISib0ihmTob8yPFNF1eQAJoRXWxklmJhUkDSPF+LH4Hoaxjsi
mv2LZoBX2k1QiDdm3ZfWngrDPq8fXJL9QHKUui21SVuDCw65vaM4PcLnwCtuGzyP
MUirdu+Gs5+oo58fg94qzmrwMhXnz8j1xnKuDwgjdCfcpXzz0udZMz3i3Y2GxKeA
eYhARXDhoE4AOPAFCKmLCzeSHX/6/N3phfLfmLuOYcvnanTOZoipnJ3M/X9e2RIR
zuY1JuIj93DShPnW9oCg5/zdpqpfZ3MBpERFgPkREH/HTCdDwwrIiStHPXDDws8d
vbmkWL799y2W0HyMxMkAwkcJGjKXjzHX4w1zXFPDvshL18VFoE0rgVgh/IIk6RY/
7CjVaqpTT04Ud/S5JznVbf/DwEAjnf6ZUWYNxu/2MxjV+qKGT3AKV+9fnB+mb00A
ICevvuzG2RaBZQyFktMoS0kbkRL6JJ8fiHDZIbBHdEh+lHhFm6DZlK1faoI28zf6
XzWI9CaZOvfMiUso3Dd7yuRoW9WyphDNNQ0BFWixCoaDd8V3zKoCUoUpsWxkqnoC
7RbM/6hqyUTLeKQYwyB8vxm5hJCbuiy9M7U9hBZE6HzxeYznEimdJPE3t7l6LVhb
rDzL/Iyqb6nMmXC5QGQAi2pMVzdul9WdP9RR+dBnrG7I+A8KAIxRRsxVwTk0iZ7F
bzffJHIcLfy6BbHjUqkN94dC0wkW+B4xZ66eqyAgWlO45+Q+njGNX0IYG+6AucCQ
bGVfPin0pIfFJemJ/7Ki5aFQ1L60xdY26eqNmGns0wAvfXd8KN83LYZV7tmTZ4BS
ojH+qZPPPOXokLmBHYBYrzz1CDcVo4uJVAsB/62cS+0ozW8PMSTQ2TXXxxdxOvd0
Kv3ahowbs04jePlC5qUygPDaeMoHs+mLTXFntWIvJ1jDF4256NkZ1oVMosBUQfHX
Nx3QkfYzhjG0tmZE9ReaOPFwLnYkjTJaSltQ0bCkVMpG6gpDczeZ3G/V903BTaEj
IhyauSRjjpFxRU4RJzWR6payH0anLpuEO4bQT+6zrAxBs0mSEhzQdwocJ8ubRS8B
5EOkXOw1Fq131SYQUVCgBCXe6PZ282llujkKDVpxQ3BoM3sOZ0psUl/UiOdhTqm6
mIDhsaX2a7YP4LeSZit5qtR7D3Vk9ZgkrpCRSQQmnOHsvCSjKGPcECuoD9FeK20B
bQuoH2anEYB7400BVBT9TF6mGkbp1JEn7houB6R8Us7xIWCWjxHnXbS8MAZUjdt/
4uSAwVsSmORCk71IZQ6sj+J11Ub9sSRHvuGMLFcrkzlePq4Wyba7JooyOiAcDtDY
GATT22DHe2tREQtiSCgzeU6sW6j9+WyZTvu0DDufD20lT0hcmgtW8lOqru7n9nGq
dV1swlqcBjXE3onKWdWTvxU6b9i5jAdJia6hffbowHHrlmRoQo/WHQR3oZjUg3c4
K53ssyU5kR7p4CG1yaIP9NgAZM/gpnKgDg+pM4a2vC7WbqD+2Edq89I3lM0JciPU
07Es0NgDigurdyjNR7YWvTDREpQ+uMwNxBRvMUZ2jxJUaxkH/68RpYqz/+mtboVI
IvOJwQnn8pNUlw8GCHGaFHw0I4kxHOpdZuu6nm/FmkyH2WQs6j9yYC0C2KYO5fpR
CompLDL5M7S6PrJsnEBQTVP9TqQV7E/YuETa+YLvWP1IwQnv5TRzLHFviiKTfAb5
kQ2115crrXDtGqlbhjPFeguR9H24EUy8TQd5jmE2VA34VMBJvMDot2ohDbNiG9+9
Ndvqi9RpCJOkSOCJHfi0lYgSuGdawBz5qGJt897vsLGZcR8DpvcFjWchjuRulLCQ
0ZB5Mc/9IxTriVT9UdNk0tuDw3VlJgpH5yVATfNWgehcZ2PAnPwwG2c8OtkU6jxa
XztBBtMAdf2Aa5UJjBeeu7uTBe8YslzIgjm8lErAuN0MdV5JurupQPrVEYYmFw7h
l9QWMqXBFCel5Kva4hPzoDZWOG7jEPnze0tNL1k4aBtp1pkC0O0vNMtGHB61/4El
SsrbZeON5eDhaFjGGpVEJjLqR9wecg6vaGZGJ1GSODzjXyg3CcVVLGdePlw7Kc+o
J10hzfflwTFRFjDowMTwqkNx4qFsIjeQGFb43Me1m54QzWDPQIE5J77yn7XzQsP9
5bthiserfmto2afoz/Er3gLcbCkdO7how0KcGrRQZnT//u3Q/4Q/qzIlaXcA7+pp
rdX2SQAPKFpXKriKouMN4LnxE9GAt2661tsPDF/rLRYFxvRGIIbZSjO9D/zNQanK
OuPvx8cRVQNJ3um8o6v3rTvuhFnCZjLlkPhAzAGBTxxFKFATbTdLcmvK9Q54vTl2
8lQGMrbsNBA6rUD/2jGl41lgazun4NrrupfmFlEQd6tIrcGqUYzafg/O7YE4ATWp
XAUco3VLl1MBAqZ7/JyT9NNV+GxhpiuaKySFi16vc3AqVVsU7N+R+IVA/JeZBlPK
D7bUOHWc3YxGlxTVX73bfZf7+4lZIQSwZJIRwZiNhay16yRe2Z50xR9NJIVteHnr
ChyAKhZRdcMSqo9aNDAlr6nzlDw4oYvFChEohlEZDn5YGfT8NPnPTV5wbk9gCYZo
jorGXqR5fiLYTbkAsHkfXL1rRf5/+tkLnVkjxBAUxLxjZscJi+j3AiTKMccegmyR
NVNz+W7LIHHI5b+lkVsOFhwT3Ibq15THptj4BL7IJm7meNOUEtBVjmaSylV098pS
oq3m9R2jXIGI0GA6uLhZtya+StMMCtRLftIcrA91WG5t4ppUS/FO/mKVv2oh1hDu
mqEDOtszBSv4yWNudqaG8MUyzP4wCDz2sIRptX07dCSlrYGRmy1JKGevr7DAZXGx
5Ogn3Ae+kTVc/CQMdTG3t9D2aVY3zzOYz/RBA6/gYVkxkgDPkjLz5nreXCQJ+dmy
+0Y3yyyZ5ZLCmYvxmc5pktLqqIzvGMgaYO7wEIc9cHlf/sqSxwWePWJkKZCTwbH4
H9zBj3F+kWuovKOhtBU74NugxlYKPYjKtvsvX3q35ssk5hQzvSnK2SmK77/uRsKL
WH4oZeMKgH7dAje8cUuWA9lIfup5xok3WTQADFTIFwrdoB3112LTB1PwmkPCyL8l
HbdtK0vyljT22OSVDuRCgXUfWhxqj9FzODt8wnIyVmq2ZMQaroujczFtelTkovpN
3ADPdajJbNvbvEaLIq+Q4NYOfQsIWA/01IilbRp+bBskoIwqQz++3Ibo04ZsvNzu
wPzM6iumIfxMAc6xOviUqQyScN61EXgR1sxVK8p+cBRQFmVge9leAQnAi/rX072T
Mp85izefB2XIrK6kwvwP7QmFacDU/aZ7UndP+lvVPuZY5NR/Q9wko0cxGa3WFAaL
Lq+N1gi2hsaTg7+FNjnGLGb/00pOxoh4OuUh0Ryswrj9++6BuB5QOy5g2FH0rOIw
I2FEk5DHDpaBgJ6H2Ay4gOjO11dHCp0fBegzlrfGT2EtlS+npcRzckrKqxg7oM2D
rab6waz0XInndSX/pGM6zcz04oH+MetapKXXhNkB9YLRYXX/Y7VxNWM7jo2wsnca
hxZi8/xzdvhZAK6LRdcLnk1b+t6DLhDwOwPWn+JlHXNOT0SAJzw39r17a0PyJL/G
2xrZrWJg+JJJLL/yWMGWgJkuzmXilRH6vWmcCT6z7lUSj9ZKMyZPY60blzLXwBJC
hrL7AXacOeKjg9jzElA4ay4vyFQdp/Hz+3xs8wpROrAequOkfyZGtc81wEPfzq+/
bnxLrvQPwyNSfJFWkyCGgBysLon2A5g8eboCP75Tth7JwP9mwBmH/w0iOKkxfmbc
tQvhzllRa8JBY7YBFkRGgbGQt2lZiaAZXAw1kbx0axdFkMj4TqsNq04Czc0D+QoM
x04RgG9G0FRw3oXP1LB49BPgW7VynzWoDw5AlcxhHbx5sXExJe8Ni25b5Q+Sj/xZ
Rop4+B5+NQ1e99osYOwN3YrGQHjn3SDeytdIG35wCdWqrpvlYoKU9LpGY5F/pGwr
FtRUxUrLnpucRk9OiLRMwRJHVMXk3jUSxB3cPRCfy2otkzw7N2kxqf/92pHho4jc
ruKlf+Cv5MF1SEfzYy9kDTP//tYVVl0I1LVQavC7vbMbSjVFaiZm3l4byFhPW2Xi
/hVz1mTGPuGriPvesB460JKJ7vXLp9a7kiaI7r47uxLYvitM3Z3EZmXT6BwiWp9b
Qsgs9dwakl1Gu+N64JRq/8iXqTMefdtuCNsAzJABoFRmc0hgVc1ZosvMVu6LdWT+
e1ZYk8jsD3+p9RVL7YW5yvwFy5oKFzwDvHMWB6aT3FDypTE7B0UiUwrJlliEvypo
J/9RmtXFdKQ+meHFwG6vE5DgHGRuAGeCWNoD6NvXYr0jbvpMSeqqfLNjyWzn1PxG
tw0oXB5MLuQEbz7Q/w/+vrO7FiZclY5HEEQsVdp5++rUJXV8Zm4OracmfiJ8roDK
cTdSNibuyQMZzF+o9E26F1DKfKhCRfvin6h/87zJr2Gq0jQJQ8IWKfYxhD+32939
wPUMPauPT5dDlzEhExWEXnwgnQnbPUr21tWLzci+ipvF6rPLx0egrJqWbmrcevzL
1rxEQUjANPa1bE69lhUi77wyv47L9I6Bk39faG0JZKVG+yEVx3KhvqIQ2tShllMq
7QEaZJBD4UQQSeuFqyxF0GU9J1Hb+rEq8Ed0t5Gcz/afmVDBbohW+uLZtfAFTtQw
XxTwPjBt1xxBzW1vC6l4/xBeCsv9vzIHB1kC22NaHCdA20VUCb7Yq3Hk9blVoSJ2
/lmqRUEnEsC/Ff6yIQn6c0iz9Ocpjx22+ZYtcnTMgVwhHt9XpaXfw5gnIQbuJJGE
q/ciqPgos6wZ7mrWxqo0N6D8BkK4pRaRWaxcXoo73HL972kpxuEkXFnBB6x/Jr/4
mNHswJNbyK0/Zzme704pBh2gr6UxHwuwQ3v2QcrQg7GGyV5DRFpYRepy3qbdcqLl
MYE3Kr2a6ZPFsSwCSMSYyMvh5wN+yaEeORome8iBrnB/Cq4vdnCzWUvOnXo6wwcA
3Zqn0/DmPoMY4CFZsEcH590hmNTAnSk9eenY61jF2LAd+lc/07YPmGk70v7oVCGu
SFmgFQzmRn1+yG8L4SdAeiVCZZPg+lLsnYi9BiF34tb6FsbILGiY2lUMH81jKi62
jEU7XUNf9XeHGDOI4g5DyXhEYKYuzSoH6cYw1BqVq5ByUZAEFz75uxnVckW8gTHo
8ZdtKqscCS6DiwGuMwAfZdWxBgYWLpTv16bVg100cllgy9iiGww9PSTzAgyiSfCM
olQ74G6EXbUugSaffG9GRIBAdpnt2yI6/ILPidwFXlIEPZ0LTsgmL6BxLDkna4RW
2lkmNdY9tfzks2pMHF0j3WddhHhHUL3ZGabKj4+YocLq0kCGzXrn06D/QT7El2Ub
eYvEDHeVNs1rbY5I6+i+qHgiMEvmEvD2qrYbOmJJ4tX0JAeSui5oEKXVEJu9w8kC
bJJXO/ornqM9Y2h0+UrP+QzYn4fw5rQ+Dh6alVHr9wb8zCXd//jKwHUowciDJvkd
/O5UYp/2y/8c0idOpyO6EOxi0vlRLt2jSTycvaLzfAoLgVkK8o3qLhpCpFUt29rX
nJt8urNh1SUxuKmtW5HPj76FPnX4rotbCtnbm7etfTFdu5DAJ/JAHNWHZUuhF6Jr
cUjZq/scGGjqRf0pHDvUJ30U70YIsxBZjXR/EzHBSUGrXYBz7FH27l2xWyviuI4k
an7VOcVfiEDSK9in0tOEEEvZEJ90b7svnFGlPlv9dlYTwOGR4+zt4MPsnPrYPbCV
N4wX4FKDonY+W6kEgUZ2OtQ3DZ9sHAKcEZzC0FXYihfmGHJI41DAEvt5oLuTDyHq
rd0IHv9ura3IneOkFb7+gNPOr+2FSHFnYW2Gg4WoZTDN0yxDxrVHgnNUm7c5BNEO
qcMfkUjccB6VR0M0gxphJj6r71TGDuMvT61ZP939KLqV3ZBYK6LUQqQoT4FMke89
irdL/xtdDjihmWTcV9MLGGAN2qLdZpHOOxOBHGddr4MnRC02Gw1eCPrh8sGSmZ57
FpldvlPWCIUSyl5Q1mbT3W8VUBdb7lMR/YW7GGevOD3F9RXfssYiVJB9QbqGUUHu
TcSU2Xq5ycn0YmWv6RuObn5EO36r5GCvAf2+H7Y4Q/6WlnnJ4Te4NGeDQQInnTxZ
MoT65DXB1PbZ74XBJdU8/m7UQBFD25mtRBKXAfjyGOb0WSfvyufJxGTU0m75RpbB
ZsUQEL4V61AcHtydWuhEswpLhAXKDiP+aGIATTyAxHm9A1MoaVSCmxRI4aO3sVPQ
yqF33Yr3ACMCSwnTARguxsdOuUjxD0Tc8ZcIDw0WtD9c8mh8XmcdhfIVNPo85zSS
iSs7Uiq5EuZcO0D4lGO8RyVy2qE8UjaXB965z9VWmhyZVIDaJO3PMxxZmdxbHMEo
nEKo7xe0YkkY0Sf0YrnmePvMH4THsjEQgQn509w1DP/SXDDUHL6UiXzaXHL5cX6p
JNRXme4ebju22rRzEJNFQ1xgRZzkfzsfhHkzG0A5cSm+FDLCiXau8toA2iyCY4qG
astUm2s5wYoG60k3noQ/mK+ieu9oIS/9A+nTIuIYNRJ2jDRoAisK0XHHoZT70PMW
g1pm7fK20H5mBQY2kP9BAA6GZOrBWQkjcInynM7mtZR9FK+Ci/ugLRq1AJ0xLNzu
Q71T+eg++WF5FKvWqABQm7G1Oy6pZngVcFu5Ze8yLw0RArK3xlkXaywRbYvjtbh/
OCAW1NzoaP1T35AW8s3EjspS6rFCAZRLxSQlL/lBANGtEfpG40hR7cy6vl8gIxwp
jL/RpJJbJJ31MEMXZaaDny80b9Ohk/NSiErDjpVoHP5jTJRBO6+p51esqFY6qHUq
cHC6gYrQryyQeMWKD/B14mgiZdFjtqDSi9Ed5EdAza+0as1pjCjMlK30HGq6QOPF
JfX4L69cf3qwyShp9YUxNf6j2XSVDppY8f7Y5ZAwW3HtzoPH18AOCC8HpXjuJKpG
/CvxAaOdVY+V26go2f7dVIDw13jSl5kYubGWpp3WbQrbFYL2E0zHVmnyucrOdMgu
pcmoKK8ZggkqamfYm8dY5yhujKkXSN0As220ts32HWzTu4f1JOam2n5o2PpbEpxr
LoD7CgJbHGEcVtoSA7nSor0yA10Af0CmsjEYL+W8lgYEMERcuDYcJKyRd3OE4f6B
+A4DdAkJNhy/X1zkyBDz/pnuXUTo31/KTYZ+dzSnrYbUHqA6FuRPt3877JCNNxVw
S/f+nNYkYQlEaf04FTfHSOuLA+WCxhpRYCilJet6tLKMeu4gUhfpICNE0rtNNoub
2qRhF4tNq3AFmRuTanI7FSOsoZb5hyKpelszGAVxeDM99bm56GVZ3LarV2XkPD6G
+LtzsnIIFrhQ2rZmCXjn7QpONvx4OLf/lnEfqxXbIPFlzM4xe557t39j7E3CZN4T
VWcUHqpXa8H0f6nNtjsPbJBFyLTq4jUPueAFLupFof82wr2HmAbfSFnCZ3+7LDXs
1+WOnr6My6kNd9Hoa9OArtgdpKHsCVmaND85dCoM+uyuTld8kVcklJKv2RT3uY9/
KAdRPNAVIVQgw1ib/6cDADuBBtOpIa7jsJNZCSQhCV/40LMFQ7HmtFRoOUDy21bq
+2liX2sQskmmrjQvOjTbAqCXGIFYY1UMU6/+j1CC2fOAxTu63zOX255KmWbGwNmQ
JMISCk69JAAp4ShdqN35i8c/c5OWOregf7Gtbu6kmxx7XJ1kVSF4hdikldHvzBJh
ayApLnlj/a3gRexUSgJKTale5cDcWbuetrt6WY5TDBh1nWNOXAYR+YhNQGlMI/J3
Yaw2aUM9GS9uzPv86VWmKN+Gpkz/ACqITqgVUoodAXLYUY8SNbCfIeTOwA28BO0f
7kDfU6Ew1xKjl8tNicFuomuYxnxr7ioi4XEvbaq08Xd5Vjr3u5rVw1z9B5DLoxOI
5PLOGaaYmkgQN6vvG+ZbctmK4/InkHued/ukEGSPkgCaRk3PsVbwHY0u/cyGzNgC
QKhabGF327C1NI0jkL3o3n4KcRODLsx/e8Vgx6qNnQ9HVYyqn5LPlwu4l9G+z9Ou
qKbLC84OA+04+F3J0OFFrJtbR/k7Nj7rnWt7EUcqImB55eBgeHdBFED62rB5GVfd
EkUr+CytNYJD2Wk+4+tknd7G4R8VxLPG3V5oHKBJM3wPmjoKcCNJg9FeyN8Qvjs7
KOtFYubpmnkIX1IEhQH4MYc9ezpAKhmy7t36WH9UmDCrITn6fyGMsU0k21uvAVdg
w+Z72f8kN1BxM9xFEvTlyZHiLUguwmgn3NHlr5vLX5+YwXbXygTjR5/P6qXg/9Rr
fIbJW/yD6TXTA/YUpLxSaEQVrjiarzQVplHldDwXdTmZxPEUquaV8N5544g32Q1f
lQSM7m2RzNEwz6JZu7WJOStxP/cNYPxgpe9zpi9hY+aUdVdY9apF8UVgXafuDwmF
qTGEv4I6ho/SinlpCweqNGmK4uPrv6SDyGPD5p1T8j4xQjZMuy+SdQKOIKsjKg58
b3AiusleoYbbkTMGWAm0euGrVh3Ym/kvrSzwvGbF1I/HwpcI7o7MV4S46Lywlmkx
izK5zVpX0CO+1/83WRz0i6EX7GrUjbqtT436vFaLwP6q5WV02HA5InecNIdJE6/X
6QCJYfAcQ4+Hozh150hDt63YwkvSjw9rcuWMYOJUXqjRSre5NSviOIpOgcZPMGuy
5xhnJg7bgC0MWWX4yslgQCiti2OmfD8FpoozYIJUnVZaaXECzgK8W/i22MCAEUj7
hTl3XIe5AystB8Q8Y4aY/tGvPRF+s+wifWgyN5tmCEB2jeWu+qyXAUCX8RyuvKL7
7XTUB6bINN34vB0i8u7p+TXWYW2kcVfucS9dBEkhCB2OBfXtwRC1kUa1ETAugHS4
KQQeDKx46eNV8G4ln0I07EM2vecZLPhjmLWz5CB1Hl4iSaLxKeRjwUnXQ+0z6fHo
CBfEmTD2ESBG3jatSKvbue6CucbrMe0/PsHwibSTcZGIsUJ/fxMNMq3QQU9jzxpc
HivrZ6UJYdB2HIIYfN8zOijsXX3J1+e6WUPWwmSq6VZs++OHqOIfQ3ihf7G6S345
2ETEVd47qc3ztoEy0JKmpwfqKUlstACcUVn5FHbm/02j3hiQQiItihbLhhkecyhC
LFkGWYq+SgNS8ztVkp9rwKtVdtmxrqhcki/cOHwFbLDJE+I5ivPIX/vbHu0NmHQB
xUNO+V1MGOS4G/pJS8JtqiChY3MpLigrXKl1ITXSo4ucApX0mvE+RFzBMYzcZE8p
YnbWBP+mcwwp5hgMh55FlN9bdRU0Yu1gFDPCULp8cIKb2u8c9UtWVrz41FVYmQMA
mqlJSutMRDvgRuFMs+sEGDJHHjUche+KGoHZD5T0GBNtoqpSgl2fyr6h+ORj6QG3
tbaCJZcwP2We5TnBfWoP8YZMAtSZYgIciac8WzQetiLvtvwOXYQCohH8BjxL/y3C
/LDIqzC0DTkr+93nICrsLb293GzFLFkHP2d5pVzEzrB/TWBcuq+3wfsyLAyJvb0E
E6ryvDZ0+pYm3J2SiwWouE8f+XVxSi+vLuy5z44kcxvzwelK9ubdQElcHlKm7hFy
2NZxLqMtKfVIcvjXTcvgPEWXBM9lDug6uIySCiowX/TXm2VY0MaGBU12zQOiyWli
ljGyRx1JiozgoVFfoXMAphNjZOU/lVU/zSTvHSksV2JdN9ubGddK8L4B7/ycAggt
MNQqIaHRROY64bB0zNKTO2LvC4cQpB4etXX7XGxuwmQMsV8z96lMEFg21y+0cMdY
PSPq7N4fVYRHDtWXPBgxG+1sWREfy96/r5sn9L/KjsREAQJbi3P9QwOk78dy+lhJ
hmhpCSK/aI0ppQd9COPimYFqv6HWaZUFWDhlPmDJoCC7usPETWwd6ztZHreDJrCk
/it1JjlUfKdVAH43O371T2j2LLaYbLnOkBXNtddtvSXJQP5X8heVUedPqjQM8cr8
3Oz8L8XS71Gs8xZVVW3ggWIKThXZnRMn/aaZFAX/5ImZYDY74qz/NEPS7y7R5tA4
e6kpQVydyMG9IPIqg+fMdhQZL0r4gJtaSHZtG1xnJYTe/XgG7I483fQzR77xsN2i
NUs/O0sAF0JrZyLxXpoNQngvHAMy6TfWWo9uYJC3fviT0yvwAeF78XrPnltip5ol
1LyevKcgwpX0O673W7aCEc96Lmdd2uiujwpJQ2CSCAaiTtR59iu9nLfhPQT9/6AO
N/ox+LZj7nmt/hSgk3EnH44+7+AnUikqhcxR4MREovQ6cemadC5plrQUfBi6+f0Y
36XZJP4xhwH8x2rYnsvm49DGYehoorrEhYBdRZtgB6ayvDk114ISjsabHxeiilw3
iVQu9BZU6oM0yuBTtwKVQ4XoYDzWAgpQjM6KRe5YTV94J5DuwTUj9LxX3g8wxOkj
6ihttZopwYs3ZrZbVHZiQkcHTZIECdjAkNCpYA6Tp6n/srUyU6OaakEhAF76nMaB
q3f/3zptQNcUJmg2NSbRFmHPlwJOQ8K3ryDoUZM/eH5/n/ehOG/GnZpvFX/V/lRF
6LDIXNqJCx1XnRZxsWKncqe/RpucC3FK/R7u6LAdo0z3uc4l9A+GG7LQFdV7kMR9
V8tRRXl+zxXX0fyFCjnCBCKqqfhRNEp083+stxd3jEnoWNxyH7grIaz0qesLFnIp
ulW5QuLCssFB5iaOEeXanNCIrkcTASff1vnbwpfz206w6+E74ycQUR48QAhKux1j
5JhkdAr25cZyGV92TjqI/OKlvWpFnGT8gZ2gEYjVBNhBav/tmVT5UVOGyRC1AAOx
Q/Gx6Z4OPnnc0egqhc+QRlFG+SfXV9kHhhX3X8h8zI/2gQQH9on3Gp9My1QkYaxk
Lc7HgF9neiKEnXuMAn4AIN+XYY8Csv153sOmwVaSTOAmy+YeJ8nBUeteBOM/qHEs
LLOBC9WX3sEPKhe7d/4r8cec7BucD8Qs8q8DO1i9puC624/Jt0WhKRSAdxwgVhDB
hwDV5szr0gvoPyifFHpXlVasrVQIdKoZdz+vNvYhkHR2mRmmFM2ZLnErlagSPkRe
9DmBEOPP5o95W8iFyreds6mOguH6N1cCfzns1hXisa3YUcfaOR5ghzD4d3mpI7ji
nnyh3d0XGXH8E/xQKM8AW3uVyO+LaLayCSWU0fHzGRkLhnEf5P4XWyHsSzT9+2R2
Op/WY6YdzswYrBMEsp7x7qIXxnJPCrJ5dUCzVYILeJHuVUfbUqdFCUJ2GnMPs25R
554gut/688W5b9OGSYLNZTtspzsQRdC/yqJhpfKR5iRlR4bG1Nxrb7ZNV7nu78Zc
9OUsSBarXqyASsgmJMN6o2zIYrZE6fztf88SiiLPwu/qNLZoOl7Yrhp3E+60pAx2
YX/pSpOlr4lLdBog0pRXp2FLeJ5s4k48CtQaCoru0CDrkj4nAK0WJMWM8bFGx42u
HOvmzXm/pooE/yU1LGMvjmGNQWaiJw4I8UvieOtqjl0KMUNwxnoqL3PCchL/XyTf
DgXfTMjTOQ6iEvEpWulmvRu10pkodFeleiwNIz5hEcRfwB/T6gLUTTqcvETaLnrQ
JJu3OZpEei154zv6V1C9jZfuHmcnzXn7zOafbjP8aRgVzSg6MI2Y80VU8dgtaivZ
M11lRfhllCIYi2ySuH2yVOjQU59+94HMfkCPCsNL8DxHC6w5iwCzUK/fvHhb6MdQ
AU8JQHY5EbOV+QGVbXWsId8+ywPHB0eMlYlc7gTYKiP3kux2Ssn5RkBG8ca2JXMH
wPvaBROh/PGiaYbvvoUu0fDem9ylSHbZF/m/Hi58zRu6q3P4gLUP7Pxvt0IOSc2d
lkJy1Tk5f8GACiXLE9EJPe+3po9WshsZTp5BV0raU85SiUPFxy4eVJk02UrYnm8h
6n8byhOBDKP6uNQGZxePHBB9viVcEbqGFCkD7rTPsS5vKlZk3dV0wPrmXbYLAE48
ETozRdyxd9Q1kZcOSo/thHebRY2rh/3UsPA/6qX5m+/dHo+zCz1gpyyXm/poMTdl
RH+/fsDqa7ajIXh2tmlLy95//z/xgfir3KenBDozsM9SNf71T6gsirK4Eel/3NAa
msYfotiAizlnlmQe4Gshm3hpWX37WrTpjlGVJarJa+3mbom7UhStSVMQBPIY0r6f
SOIEdoYoFJgIaErAy2vJRmqRqea+Vhg6o9nPqXveys73Ls5mi3wGY9LgvUCF4wcp
X8mlNQ0Xa0MUHWx7/K6sww9UgHAXOj7AAmriipagjq3vzZb/4iBYh3MDZAEbdTJE
nV9hk9DxJpk0cNwxeIn7VFLixGZGNnDXyPTSjEg7qYiODWHTDlAFmeU2TaOiwOxv
ZBRe9iQP8LAKW4vUwGaV2YcheXmg+a3VhTslFlC6Mow1SGjo3CQf4hddGAUbWXnR
2rfwYI+OSBxHcv4YMf2zhDaOgywNhM7+ennQDKb9h6ysqSfgI1tVpn3oAhTwhxgT
LRVAgPNn4+q724Z3BYBx5fuQqBlWr9gXM15D1HjoNxIBRqrhAdflBpNlQx2T+lQi
iwL/mw5Tm43P/sn+9fpRJFRENQlv2bC3R82T/t/pk0BLEBRU46Ilt2Ppb+oU5Jzd
ANfo6Yz7j9AiJkmj27B9tTRAuoK6lRu4GR3a+tB+mUukkLtAUALO8vKVqof9h0dG
ZEkRVy0OEmhmq8EqZEEnbmKA/FyV6z60zm89ipKZ4x4iGalfayW5QDYxX2/2Zm3e
dMuKXjTpIRRCcUwVs8I8ZhbLTl0vFRt34kX6f9Yd86hEge374UngB3qBqXWb8emq
lfbUa7Pt7Oxp4o0LuCJEDEuqjNBF0IOKjyXub1z+UbxJcoiyVqwtGb1F1vn6sQ1q
a0wuSujrR+HOZKRgwRJ5G+GY8FWiJ/CUh8+3QLhawnoSEiyUIHMEqvCkEy+FClVG
4hhvMCb7RpS174myAMzz4mHV46MvOn/crTvWk3yjSvOB7Qcet0MWDKJUNISG39qu
/AVEskXgT6I6jLWdhQ17ycSg0Zc8DXZaKk/+oZrjY35Q42dMrRotJTpTIabp2hCb
wRimhoqU9yNCPP1FuFarqSysT5zVt29XEbDgWyM+ha4JTlhfBBz5Nsxnjx53OhzT
dE9VomMcxB9uGBSdYm5Ku8YLapmpwIQWtZBUgV6c/MVGmSuMprDZzacaGWknaM5t
rCZdrWelor9ARf3SEEN4R+2tAyZNB9HRASjCCYcs7q8oetHIvZLaqsCCWrVPsM4W
6OC7tHttAxuW9Ky5OoJvs5B97e9B1/K4hVn45+4/6JuRsv2BPMi5ka0tggLYkvU2
7C3QLTOh3N3NfHlrjHv35GBYwOHTdMV4/WS/l/1L/vy/xLgMZvfeGeT6sTyOSPMT
X3ySJ//iPtnl2FBWFS2JhG9ucUoXH9CT003l5D+kBLLjgv78dtZyl/NNpOPT5OQ6
2X61OGbnCJ01TguT9z4yG6VwiachAkG9uiQRjD7V4dfCSre9yBloS+fYvqmdXr/I
vJkOcULMEdhIAS2DzDy4C7PPidrhZaRU/aq+NylgkvIZSKL892grA2ZW8sa04/Qx
ndVeGLD6xr2aWw0UZJZ3m1QB7VMPS7Q0ME7Wb1hCsgU0pL1bE/2mNWw8yhrcK7jn
3zNxAWBrCta+qjgbE5+vWALLcDh32ad0AVqXpkmL7faPnNXSzdDbXSbQm+xzrpJd
URJK0lf3IbsBr9ZeI6JVNmyqB9uMXrJ0IVxsa1fmt/c002TeLHHiLjznsMG34gYX
6uPJyyOaftMPXBxIbDrLSOg+Ai2p5CjJa1d96H/5Sr0XbfXOTeYfaxsiligAhLzo
qfjuq1ljTwZDdnAe3U1aprGKmug6w3MwUgNpYcPFwkhffuFp5PfU4WOLOfX12eNQ
lC7d7YIEJtvAQMoueOsAQ6QvHyDCd88YO3YEnwWOZYfXlvbfmMKVudKGD5zIWwJG
0oBxAkbsQIyUttu9q1Kcsv6e+I9+esTBSkfyeS6OWYSW/a8POX1TPw9qLvh2HbOT
V6GD1Y/iLwx/8Bj2tpuJAaipY1s4u/B47+SQgEI0djFsnQr7T4jRooI/xC3tF29K
4pH2m1KRGT/7S6namn5gS9eN5HnJTXLhVI5EMWpyXZvdk2qBdmrl7VrSdGpj2bKl
YbOEFOTYBVZY8klyfZnfZEfs0ZES2lm0539G0pyW6wBQ7IWETMsPnH6/mMkFZi7i
HNpCrFAMH2RgM+7lOPZMnFXNkNH/7b5pso8w2M7GWuu40x1blsZf+WIHx5KS+t/P
upV3RiuVEzKVebDKIgF1rXbQllKA7f/tlwKz06zb2c6Yjb4/pltTrsOyt141o+ca
1CIFDxueiIasZYiv0zkSfSkJQhANCptYc7wTG6WfLT+9JSRPeBseFPSbVDXiHs6R
JC5FhLqR4OBmOBJ2QR11trCdKBFnGvIulKQ/9ydwwxO/kC4BhYc7t5GZquNWHNI7
PSyiexHjB/O3R0QJfi1dcs3bDRQrbKbcjH/HzsBvepmZtbHxOaQxQaYTw1nIMb/i
QTYPYYIJMM/k5DTkEZo4559GFG1c2GA4/nlHIsfo3My+SGANne5ZjzhAhy4mZ9Wi
/cEnfkw0L4xks2jVltfLu9J+yzbKHg5FUPZnwEX0mT9bYL43Hlc12NQpIPynv7Vi
IK3rFjqkfLQcow4yDYq4uYOHZfuCADngE/xb0RV7dK5mo6bCzcKwpDnRrFHRJtUZ
UG45QuQd2TBzdsx7CzB+ZgksB/xD0YKw4GL8NKhZv2+CJsA9tqi3RSThBOTkXCi+
gswrvurEkW0XFOO3RdYaPXASKa/T+jh1xjmpRy+ADo1EJrUechXUcG9pQSOxPAKc
hSel4OaefxPJv2r9szr06aLBUFTGHenTsApFEtabEGkb22QFMOzMuNZ7kFeS09Rm
q57bDOR3ICzm4IazwnQuONfwGJP/H7R0we/zSC16BVaf0eJM7puc7omVSeWQHBQK
1tOcN41RkPdy4rXdtN9npndAknxTT0sR20P5BBQ+/qEZXjPwPlb8xXqf8L5WNoKM
OipWQpEGFxP0OrJC1vG4ljmXASZkQPWljsWTzKcoXzPKCPN1fICuRAZxYimmryD9
6c4nxukOL2hqNQeAmT0xIU6URd/WF7pPkGLDChXC8bRcrOVxRT0SUQ6EgrK+di9U
D7kDUqJrnpGgAn8lStZUUAf1nutKIs4Xxqv8mvjxLq2FyxOZlrinaqj0494M+Get
APqkVRfXMMGVXh8ABUqQ4YRXTFDf0J9mNkKjvQ3IDwLZfN/M/zZOjQ7ZCfNadzqv
mM2n1HQH9y2kCzQL0RwXRQ8oFyAYALaEuW1YPY5Xt1I7pRO///i7T4UEvA0MPplI
66LdkkdZu2iN7YlmbRbJG+SauC8FnYJSI//FZpqH/DyGeJ7jnhr6VEFPxa2G4/yi
Z88e7I2+2pKP1Ox/uVbHBTa7suwuzZMHuHrPqzC/08BUugFLQ0LOQkK95mQ92CBs
mH7GfHkmKEaG3Hiwlj9XvNlRPQ1cVMygudDxTbhgv1rKSgqmlkqE6riHnjzIoywx
38J25nKtmHm8/aF46vZcXkuTx6b0dEn8TvQMtIg1c98hlLeGkfxfnM2EqAesrTSU
LKl9c+rn5l+75kixrDr0Hs4krI1b5CiiX8EFbhlubN25g+5NEjD8j4XJR3Vcq+Df
q8WxsCh7Py8QMEu99RRT8AQHwTN9xpy0ECHxSw5cHT0AhJeg+fIk7aEfxr+ME0Yb
WI8FirRtI78WTQOfHO2o7Aa6pKv5j1XG+4jaeSgB0OaNr3Pogzwvkvg1KzofNmNm
VK73sZCuS9ik/K3rUmeflHkPIwV/BJlprkvcWYZmxShYkJ4nV+KVl6AkH/8m9YH9
DNar17r7ZErXlkvrVXWp9kGcqGrVxo7GKtghAI7IMNzLfx8cTfRSM8wQGeNKlt7E
i/cvSZb3+LFW38Npm7ceucks7h83KkCwqkX/9Cmq4ygkB9OEKPN9En0i98NtCQuu
FeO9mLUMljyPSXg01cFSC25HftoHLETktpYsfleGXQB1/iK/F0ovklgCqg/yln1E
KAw62GExgUDgrWAuYxL/RNARcOW1jul6XQ5XvzukvRLM/Igl6UPavJhHoQ05IUxV
H+oV91k7yjLT3kxe+o6PjLR8qNMUD1E4LPDKvFjUdUVeffOt8OTxAc/42hw0FFba
Nda7XkATKfUHRRCkfRmOUv8UeyHiqFL1Y5ZJOZyAgNxp7RGqKifvKFdW6OfVErkC
1S+K1bt6dcgmkroB6dhWXphS6CCUbW1lrMErVHaQzOG3YngTkkwdhiKFRcqRLqKf
zhhs0wXdg/BcP2N0fOuEQYlyIz1qrPdIF8GnJKU+W4gYQQZbbVrvTHqCnap5gCLl
3nfYtANEfuuxQKH2V6tbjZPh5blo/IGIxd6dpOE6+dzLTSmHEHjzL7hncdXXN+f1
8FCOG5x8IfQ8LESyoHLlm0/XD89wb6qA32l7nV5lN0PvCPwdcIFdaEbQmUgZXa2e
iOyMRAPdCmb6ffDpA7/YxuvfhJcUhXfF8Xo48SSZAj0ZbQS9wlRLLu9hzn3TEm2c
YdG++JrxOT7Rv+r1et/j9QsrbS+/FLKkSI5Ft8qsl6ashDXwofsaA99NhTHRzWvr
0oTdVkbsl9xJGoMfa8NjOfbyOIatcxZdaUcyztJX4ol7YDFN2LVFv0VfNmQorSjG
glwbmatMRq7j3HWP0xQTZE/nAf/Y9mtv1nXIXPllPim7efhRYZPBLsrOAzrs0j3C
QDTTqDA6UQHaKUdhD4B9BowkufpHDpMwqeFpTqu6vIzjgkx92sqPDsTsU43zkr36
R0yWtMtAUxJOi1zUtW3ODeEdpdbVHpAUbtL3tO7B7L8bLSebvCkUMBrcFDAVb6Ds
e2qINCEp4Zg3JEiO3zEpS0s96OMtGood7Lv3bY3SuD6mD65JTG0NCGAahKUmIHN1
rVMv2OBxdgRiiOo7E+VokpPYo4/7vNcP3Hb2IM8H1DguThBa9nC+8qmBvKrCCD04
2eO41xwcO3pnlyru+u3Z5JGfWFCrfxwNm3EsTDH+KLVP08x4vsBPVh+ThG4coMhV
lZ1OspOn5NktiHs/QMpR4RdLp8cekQ3rCvkO9yQMuUv8EhyF43D6uIhamgCuB85E
zArAcNbEr/3XC5bQp0c+rwNtSMSd96Fgvrvlwr0vwyusrlVxYjqL0cd7bAZU3LQB
q8Y+rvc/mvNxloUcbTYosdyYu0J++md7YA+YI9j6u+fVc60HkL8wusx5EYgeC6pd
B1tU2kYPGyiDM84Ao/Qq0H/ww2KSxHvuGx3PwVCtIwdnNzydzAn6pXGupJRNOHWV
cc97b4YpojuRpj5E8quIy/rY5VjPoulMh1oMKXyXdQO5o24kSM9JOWCFfypNn4dZ
Kn1Qc0GNdKe+2euk16Na3y3mDlaciI2bFpQi7TlCufRupIOBF3BX90JrO0K8oUGv
bdbMK7nGWET/jlTdsiUbZgyhRxZjBw9O8942gluNo/BAibSPkRmYg8SbneS7AJoh
9UjHjZC7Mxg+ZZCd9cZZOwNX2c/jQwP8+88URWnWikrJvxxxrVtFEdlZXWVjIY9H
3FjQWnbbzz1vYUHb8dwvzmLvnLZpiX2I3PWmdaQsLG6M9ZuJG6/0jpslHT+YjGAv
QEhwotkEuaihfFGvx358xmupUaD2G7laUWE6SonptIVl8Ny9T2zRq61jv0IX1q/l
0uLighEZcr/cWjDO/qy2hAYNecdqcpMrpl3c/0SHkAx+cpOWIircu6H5ne6VaZ9t
dCl401FgiUh+XuHx/3JnCipGfJ0GOZOvuKFdz/kbCEodE70B2qtCpaL1aoX2gm+C
LCwrf6RjCHPHGQkLiWN+QN8gJRuuRzyP6gxgGAZU2DRZdarvsC5uBApL3Axuzs63
8Cj8mkA9kzhE9wb2RPexqoHJZHA1ov440UqUPJ1cA/CSC0PBj6CNp2AzoniarTm1
plNUNPmBuX2LxutAq+kWNZkV25fm8qD2MTvaZQa3oDXoWFylseuGMuvnoTaxFD+6
YXpCmQx1iVXoEdgR0FAfBTLS6cUrvStEmm7t8tDQMrd+kJ9PZV+Z9Lj1wYVlPjqg
CK087NZNaOpcZY+Ts7xpF1tAvInddhaio50hHi7vGnjxQLY5zOmJ09qvf9zI+sef
iBj4eWlULCNeFgRuAcuyjMjjBOGZOVeF35n6d9mHZ/FrtlBMnysXM3/gXI0tOlxz
9u0Zck/M6gQ5lhQLx++RyYIw4lczjkG3ocMJd627YCC9QHw+Ab93jefqQxwUNgDX
AKAxz16PFkc/FZHa9sv2d7ix8iIgWTaSdD3XDEIUQTYZkL9dlZ9xERHXUO3lqmYu
ouyX4dpAJV57lKD1ckyhAujxH51EEGtrc1Pz00nX2Q6r5WiYflaSyHPu4F/64e2l
VIdt3O5HXV+7Xuc4FoFoZMjU2w15dOZ3b8iNH6+6RNmQ+UmUOhUY3vfMVBBNt3OD
YOq3wKoxxw2/mkST6W2oNzQGwppfw7Z2949LrPgpOsrVqRe4ba560kjlKu8neQiG
7n4hOeubcwwEtBNI/pX+yN311pIiOKyBWdTODZel+aCm+I5IuzSOPJWhYIa88xOJ
5jxOTHkR9jMq12O20BtrBVLe9WLE0sByQYn88zefElsW1P1Ia8uUvAgeq+F1v2Jl
C1YpWJ0yhaeZNtnqJTop3Ewg7J3i2T2sx+w2CzlP2WZ7g4wHY02tDGtVubkjrEUB
ZMhDrFytpXfE2Jx7+GPV7C0m4yZdQpID+BggxfxIMkCbUtczRF29LMTrBfaCdc9Q
9h9ccaXmT6FQdxhrH7CkqHMt+3+9cw+34NvbErRQFfOiitrhU8WDBYWMBhldlA3O
GX4NCOIDbxTnA0lxf+P0/0shKKFBB3/Y7p8tZO/qSaATiNAY8hLAYOTnw/+KxjJp
behVDsi9N54iDpb4YyffH/jRrct/0b4+HU7zCMNt+lTmQtsrvDD4dzP4BzR4EQq4
VubhbUeL3/LEHavD9KGq2Sq+jhXPSA+0BdEfcjwgIeGs9zEn4gSrIDp0377Ut7tV
30G488J1hcba8zd0gcrukCiWHpP4m6HlrEoM8k4+V6zTROY94eLbSSzubcfaSTuB
ynWq4hTo7O9Gal1iWB/ABDkSAq8BmAI3seD/S1KnPC8VuyUKCoEfhcTw7FKHrrkw
1burACgZeAf1DtuyPhnIUQpCw5ReLv70PpUzghbB+Ej7SG7oZD728M9VGor9NGf1
u5blls1eoAzbc0XDt7J7rLu5PMEXCxvVCE2UHELr1vD5ia+NihdK5qf1K5hRvL79
4GNPKP7Rg/nejvAJ9CKGa76LMyRuU9I28+mzjMID5NYLCcIgnC/h3RmCnSdgdUsd
ksDQSNntzgP8byKVVMsqKWmJAW1Tv42KzW4lZyVZG4YkGnELNnkv4qTNEpZcYg9o
atAIzmrH7Qh6k8CqDP+pwgT+w1Eg3fPiGthAul8DoRPFCAnpcWALRboX2oEoh5Qb
l40m1Uqm67rm4zyHDu+/uVmkeY/NQGMc8PN+/pUlKShix8Qq/5uteTbxWfX2pqaM
8VFR5pL1CHVUITicTEP07NznHw+DQIa+5osx2gD74+rqHSKKDrhjVqo/pOMRodag
y2GCytc07Ss9egjQZ2HsMVBK1WC8esg+tpPoKVcj3KbQ745Js/GtpmopBx6NxICw
NIJtQAK+aRt/sSSRCOuQfT6kFNOe21LAaoMpjcXthIm0HP3mwyFAA+zuMyZkUT9Y
uCt8VodiQRHp34SgMucVNFfVFqHoF4m06Pppti7DlWVXoSnRsmEzBdF/o6MaeY1a
QgQYQ1y2AB8UyyXdaRaAUhV/rO8GRpzhEUUZV2mNCs7cu3bwCZy8OepyUZOciwF5
bNqQPVjR92L56gNTso6nXJmkvBsa3low9YozjxDBQiNeVF4nwyBHcATP40up546J
W6A0MW788Bcmb2L5WWXRkIGs1d5vRpO1CdbVVGE2v7/fkYxr5HVRfw50x0H8rTVE
2J9rjcfMxyN5v7tC7gK18t99iv0g/DBRWWNufzBWymC5GiEcnA7fqX36mTsRS2TH
cgnbhOMZ3jeKIapqAn2R0aYUVVzOnSnuZ+IGlkrJVSnyIWYtMUErwJ9WfjCi9Gfx
oCgP2WP7YYSJ2RzbBnVgilE7Sskd/ypItE1sNtIvu2dYVKkwKqT3QhBvSmMlFp8F
Vbpth31DTGWem/0+UEYzgGGGs2ulp+gBaX7GHgFY83FmCA1VhwhVn9SRoaku0T6/
VUjlkZgJ9FmqhzyvJptcPwvv111M8OdqXr/KGNKLZYe8IlEBnMXt3Thpups0kogK
64UWrWxZgoSWshFxOSqN/hCYaB/0rye06UdgBzlMAyIKJhG9V8JOKs2VG7QY9IWW
bRO0B9vE7LgNE73Hbdb8aqZ3D7CtkeMSQXOi2VOG4Bs/aHkbcvDDYnqAMc49hcis
iF5mvIWBJ1RkKOBdfDxs1b8IogiawCvXLz8znhput+XewjlDqRXAgViZcpVfkT/L
nop+tixtN3USB4ick+u7Ot2GN7eBcuT8EcASSDMycS9wb4nKb24Ks1LRJjJG3i4p
l6d7V3O6HmjgmfulKXNR/iodohUXLNqe3YaEhPO0cOVxEXfH0BOajOfaqV8uuzJS
jMMjzRQNsJ/q51tD/h8HO14jz9qmhjmXSrRb98ZhWr4go4kDmlezimq5eysHUA13
sJZDnbT0+5nxQcMJUrB5HvhKHExU+so16xpmokYBO9puyfXTjHD4fc191w6M6niz
2lJ8isgfR3cPLSKqKs7184XbGWTFgZKSJu+v8LM+m7rOT30TUa2QCdBf4kcG9Ei3
jj4ITDXh7nKr043OpBnhy3bwU9NiKtltB3Q7Lkfiu4LyNRH3a4g6+27qee9CwaBO
vbrqlUljtFCXGhA9JngpRjDQB7NjiiE3+D6/y8jfq685VBzgHAKHDLTRfp6zTR+G
09C+lm7nRhHD7Ia4S82kIq/4zXLRQgKFyUTOAcbFPI2JEqHeUIq1UnG+eLaXMDGa
9f9lgJ52JfeGLaUhaO/jbkNtS9Opdw9zYzfT+nu9aIU50AeFO9+NUB8vS/KeetRD
D6JWJCi+R0ROdPyBsV8ovEXFdxfizsjaKhQXpJ7T0vB1wu7QyC8exmQlp5nVlpjd
M+C3ltMht4OqO5SSv9yCW5FyBaKl1GkGhd/ZwRjd4/nx0IqvF8qHPDrkclLbcISg
VVwQBGv9j6eaoYB+F7vLma8PEOUwFVL+vYBQ1Zsaw5/5olOgq/dZ2ANErIBAYeyO
LaDyguuW+3mWq8jaHipFGr41SbIYJqbfEzII2k2tBD8EKBKLIJ89zOKrHgXVBKKv
x2bH3sOiXxB1aciooKSRtCrcSx4NYDyuinY2G33v9rGYaAczt7/Yx7OR61JPrcSs
IvPxAcnnBWoiMcAW0CMSknItB3bjMA5B+3OjlfDJQvoNnpoSUEAkYOBnl/d+HxfS
zE/6lnD8ua5Sh80ILY0W07/onNBVib794L9HyREGa1w1euYugjLUnCV8f/jhi/YG
jeqmbkY01TxJqeJ+jKUru2GEEDuBbv12OST4aLbQl44xMCxG3LtSb743cFl1CpaI
RgRf/muubOHekYqV49TTjffmximevPXeIPvaJHahjDQMEdxsO8Q2WZuxDBNw6zRf
0mC4atx2IiNrvlc6SM2MOWgbdFPgdIjzR/A33nkR8ROrnCW6gbpG8W2oeH29hD+l
Rml5W+1Db4UqaLh+THbbYj/7wRwfozkilQl+4xZRVCU4uRA0UobjWq5q8QmFSkv1
QJADzixZkQiI9g0NFhz8K38wBN9M0dIVw85t+Tniz+YrZDZL4JCbw/zw21p47RqV
WFUTt/r5nqz2u1gPoPHuj+aVPjDeLB5+MVyo+PAc9BJakth/ETEBPVfV0Q72+DUk
SEygrTKrPjc4b7WC15KY76728tqVHAuVuzSjcOqqM90M2sVacth8NaDbDenE5coY
/sjR5U0+21lh9DJSa9nXdQfIwfe/3r1l1GYMchpkqEhIkZtvoUzPuntg+InUSN5/
vOAouCkpe8D2Q9Z1rhe2npmbljsG3wr57SbGTH/vPVjrljJS23K0JMDUghT/zJSu
oHPY8kcF0JM/JRZjiG6yiiI3gxSSWrqo+OGV/+cCSgb344YPrdes+B/cAZLCxVbk
Qjnu2oXwySXu3akiS+jDrxE2uSPyaKFWug9zXzI7lwvMXyD/4DVM1M7G/Z6kT+G6
R4zvBgpsGJiVaXcQYOpqLTupPNQlF/V73pGA/ttaYvIYRY6mrIKkUkyL6JiagLM7
6hiqiM6JgSyTOoZDN2j27UEeZCLgJL2cU7nYelc8uq9n9Acm6tstDH63upiWTgDZ
LfufkHwRfSNJBYFCkEkRWy/ivuui9hrCfBcwcHsuWCTCbiQLapEcOLwHR+Cjxu9G
ZujztoS9gm/yGeyQCsuM/ihPfQD82C53oopBXn7bl1avjPRMGzXYwl5mCnY3oJZZ
vuE+eeUN8YELW2730axiaTBxmx09f+GhshXPasgI9K/PoFeTAizFAbUr1nyH8kHi
Nu2a2PDdGxNwmdgdvGr2wX01hAyGJeAzDqqNWh772B+Atxky/5uTuwnSSeCe1Qep
RFgEtwE/tsWYb1p20EHa+4BcvYcFvKbn4KA+9v9gyHLtgbFYZHz3Z2DG6qbPesfd
f97oAMAS7Ed92a7hRgxHR9xHzPeIXNn5wDR57T3z38+DBPXaL2yK/t+pCuHAYi/g
Byd1ExF8r2YoRnem/HDhUvH313A+HahYnWe0GTFHB9oVF/nWLAHHWw8j8l0wwplD
ZRxBzleBQ7wrFOh/CbK9kgVdcxUZ0VL5f7hZ7KOA0CwKsPDb/xbTNrl8YlLeb9yX
jfBpFJDrrujv43TMlJQli+fejBazxsC7zd49ULQEcyohEcQXJbE3StzTQANcI1YK
WCKKNGqFxKhJQnufY0KjyEGXeSyww9MnhUfkdCq/+ZcaZt8uJ83lrNvs0oD4Oonl
WKo+M5lZURbIovqE+joA4Q6tMWtYVNhgdTjpM1+EIdZ2SF6Yrjx+PQz7Snq4FlCn
Dj2yLakV1vpmwW8r8M5ybvazGMKm+29IH3KshbnlhMb3yRU5SBZyaixwJIv3cUsZ
EKsHgzD4DyZikXRE/+PgWcrN+AezSJKZXNGKRU0hbcs1BwoB1SQVTW1dOkOgQ1au
IEui6UDVaAhIfg+D6KoT71/yFtHVgNVO6Zkjk1oWruRycLPmGO3QxC7ifZxLg+I5
dwQdkAqmqZ6YOd22hRPO+n4rlmGrNSc2eimsMIgL5UG7468CkLLU5AtEB0JiqAex
enjj0AVH8YXpB2ttQXuPPU9sWdVzrMi4APd+L4KrHwFQj6/HltIlH36ZZnnXtVAA
SDm/CWTMXJ0fZpF9reK5Vv5xLw515OySiM3T6jncV/zzxBPzMRwDmljZ9/oc1Bxr
wEYqU4wQgEkSCWQlTmdUf5NXla1/aMsrrWTNYKRTAvrSNaKED8/hQSAltLStHZl/
GEdn8c0j2DJYiJ37Hg4DUEbGZo9GGcGTEY1tTiT/4xicHOBgIJIuuR6+XDbeqpO1
sSNTf0KZK2neBzA8GJY5ZQH0swJVqkH2U87KjrtI+aozCShlaiyzqiWC+azSywl7
cc+NAWAx4cfBIs6czHqHFkuFAUAayjfb9pNcemhYGSrohSSrBu37SsfKIO6FI2fb
jlpz4QwQpRc+PkwDCWBcrXf1Qt+6qAVokxvU/aJhr4gZ2dSXGN24fb6BAhEAhmUO
W7RbiSGeS620iE/yJ04RRCWbMb1N/gsvDu4Jt6EPS14sH1Sr3P3ZZLoQ2ktF2T/e
c4ZlTZpMkhYv90lKGKb3UlLwgzcEOQtwK3wB9vdYF1YjTXQ4LDu+YBxcuWhgnLAu
dyAMpSB231X2kyaJFVF2m+paCqONBceMYWX5nAoj0N1prO4HuN5i+Q+qZ/8BcBJq
5uuRoexyvGJkyWOBU5Us6wGczkeExy0b8NCZprbz7DZzEZXkcsb0wudCmGNL049I
FhCvFmMTYKjocOdAG87KyQo1w/rhRqkEJYP5JZdJrtWKMevdlUiqKU5tjURtJ3Wo
MzxE01HodqsUCIWG54kUU7jzlkzX2feGpUNa1DBW7D3lQUb/IwbZkEh4zLYKqZsA
4Pn8x/pctXNVMUAgVPRr0hmtlB3+Tj5PtTJJn+YhhOoJ5yA7d2up8A+fsbDYlqqc
IFry4lp1ILwdMHwzNEKKNS+2PkBQDVb2fmsZcxI0pc56YsxyW75/HHfAHZ+vzGOw
ybH334oUFjqEvAgz/5I4RnGE/CsNLbBSQ/ojk8ix6z/+2iCs6r87Nlk1b1cuedRD
fF7r1uL+26oGBX2oNAMUBCn6D64qZcAA7/WkM2ZBOeRaCFFVUt2xPwWMFGzXqhSd
XG6bEYRtemh1P4d9YnzoeIZVv0Nf+2uRqVe58cg+S6E=
`pragma protect end_protected
