// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
SD1w0Sf4LhDSAuLuglcIktKHNMiGL8A0007MrMj0nn4ffy0tqs1s1OzFlqFj8pbIFjsMDfnqtgfD
ut/NqwwBJzZs9mlH6iBh/WQa29n5Ze3Hf88U2Jf+1ltcWzWT/OIWxveW5o84a/6BWfGFfWOpuAxZ
8jY+CmdHbSDt3Bzk9zAVJYzr0S3WkhmQESjEef2P/6MLtE/eBKv+TidtXtOrYXzoglIsrNuOBjex
Qkc5IAqQr+jAAJ/L17qx36JPXgHNq4sPaISI6w71ef617CMO++u/35SUy8cx50tZUtQSyYrNGz1S
YTEDb+FtcAgYOEdPmQWTSLx0u+05vrXu840cTQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
B10WV+fUzPLGKE31Nkxq/0dku6MFqb56aSFz0UTf7aWk3XKLuWDpOnTv2tPTWIrpEOP9NJFoOk72
LgSLoQUUmUYYre8bsC4MCQcvuQZ9yoh4dGbtLLVz1XDcShh8Dssz98f56ptCp6RGpPwqvL29Vhm3
mKeBjgVpsg/zXtVbmbf1jITX01nsi1FhYzHvoJMSWrwsdJcX2kV5jTCsX/LCOWpal136vlVCcIdh
Jk++gTG9tabuglCZFFrTaMCMqEXwuZLgSMj58BnqJAYuYEy1ibGJG9aOFUJyBph63egz3kgVbOXK
YP83XxqjVQtuXHHhEOnJSQ218kkJqhmd6hP/SzjbeAbVJt/rqgVtnVEgUf5ILFluBBOBIKWxJL3y
KWeO6E1obR9I0Wq9AibIv/Bh4aFpmvZ1BROxsLmB0awZUFEDc6RyqHtjszixf+aOkvhdgGCItx22
mxzZ5vRQK4+jecNho8gfs+A3IzzjRbziiok2D9FcEjBGCkwc+pVWzqmiILA5AU8CTdabSuibQfWa
J2B4komnKvJ4/F2twa1PkRMjaHB3R5QIM9KHSopi9WPFmh41QDgYo6I1StPm+n2SeAjrX6HQeV60
aSpVQjopsjN3hmCo7AbNtV9jRA1Lx4E9xLyIW3927FUX830Gq497WkR1QE1gs/94H628Y9RTessZ
I8gT9ofmqG/vBOFpXee/K7ep+O+c8Yu3vylSHxz9l3elovxgL6GE2vyED8UjMq/gNDn+NLd25aF0
Oyuqg1eMoS2TY59Tis4olXyvmtBdPmPEgJZ/vKgvSROe04jusM9O+eK3XGte00b1z9YuWCFvxERJ
Jr8cLuPeTOW8xj0ipa5Ymv2IzvCIvvLT3umerb6/ZdUXG+kH1K9F++BxfxUcF1Ur6RoefakP8g1y
9oxafaOJ29qMsAFW45AlcJw2rSonTuigHpGXZk1kfX7zsAJ2fD2sU86kjOvz9/9c5axK0C7wELFR
Ldf2lex9brAJDSIwuTg2Z/sVKJB2hOucEPTv5FyLdAiNAINDXlxk+KjJUBOgX7aOH0kklw9kyD9z
ecPom2b7wGq76Ru5HpIoMz77vH4hZuXHDjglNiCx5ID0yFE3ULP3GhbGYWDg0iD2dzvcZdWPLgjZ
sHhKK5whddsTLgoXoC/j09ksf0XK06PpcqxYMvWOUcliQRU4STYMjONkTpBaaBtlLOGojnCYja8+
snB4pLgG9M9qWtGCllgz4KAL/JKWoxJOuqzy6rkdxKHw07GnADL8wxzjP9HxBqXijm0yf/ffjThZ
MMhD4b4cNrZt61EteGvtmphYp4OcEqxE1hvyj1sLItELZlZ1zQ+dqNfIS1TIYAFQgMjmNm9Tc5rH
X8LMCLZlfo3yXgwfQc21XXcl/yp01GfKlb/vRLLhJ0De4C57VpgtGuyutg8TDsuc56oadthM3VeE
lakxkWuz6o1kjBJQwU0JoL7cAjx7lbRbYdH7iJMU+OJ14IFM1gKtS19tISm2O9hgqTPDKNgoSJk8
J8t3zLXPfqlq11EIJxtsCsGmgeSDKQ3Os63gH20jK6C7bSFHZt1TSSP2ax/FEHjq0oC/4mEwX3gA
i12VnF2PttcMORdmoATBlC/Rk7JXB8unFb7kjFdxR7O7FXvyu8aOtigrw6uu9haIJhjOmls5EkD9
GDBH/yxRsxu8SxsrNJoV5kwkc2XgdhRNYVI9Ke5Hu1YwnhiXTwOIccHTTlUjf3HB/Ubay7NDZ9lP
kjQXcSGNc+RT0JTvIY+lC8i+9Wk1W6KDp1AwccwK0d6QMYWZwrhOEY9crEKuLbzu7ls5Ny4agxzL
KiaSgjhNNzZHazzZhFsNfgIbuJsWmjRpSByXe3elFc+bkQy2VDV6HB2aygUPCKLnjGPAE/4lx1ZM
5l1zvi9GOxnU7GCPYJzolES81FxZATom9vbhkn0PjSQylgqfl8gWqs54qLt9Hr1znKfQWrdvsMx9
S2sBxpggtVbqHC/+Vh93msgF23a63Wb4SEn0LHeLWnZ/9U4VixFDTl92A7NFfaq/sGKfZLEO7QuN
vGax7Fpu04pANA6YFK/coJJxtcPajlI8oj/f5x8vnrciVa1lW/61MifkWJ9ZZGaG+8asY8ifPnu5
CsSCjn9DXcsedB4NNAId0JmXY1CwwKEU5w3rohxvrUVWFwejymmoOGZDwxSJHvfz8953O2ar2iZF
LyrNLBxRETDFxfWw59XUYZsd6YvSvLfc8/AbUOafofxW/I3tVlqRY4DjDj2kKnNgccOF1pS4rsVH
VbtVv9mx91eiUGBo6adu2JUp+hNvVGX/BsEvlC98Csv3iux21g7Ugu44fFOc0WOLP0J4zTczVVv+
Rzgs6KlSk6mbJQcjS9x+IMQ0/JjdqopkWhSovOtC3oKm2WHz37QjET0RUGohuwdG3qQWuAGqQYe0
qtTGaIaAhz+S9kWdusd1P4zwGPNb8zYc+hHo8OwtTdFaPWYQXtKjMkc3nrS62/S6o5W3DFCCHKE2
lv9Xn4LU1+60orsMOZT3Tj7ihw1/ShBjTFRhFfSwL44cSb1xPGVEAeVN9aZ8lqywwiOM9bdpr6Q9
F2bcchAxPoSokeyYrGxmYKuCBCpuqRT8yv2Tu5NVBr0UxD/VgcR1QPYsHCn9Pw0TkxBTKtVtDceL
L7mWtQpPB7HD5U363fFjEyy5MX9k1WDri5HC7F3jt3/FraTJU11SkQy+2SmDGPHsUHkiVtKQW0FM
GPKjfVldJ/NRGW4ZexDWMTuCpYXe6kKuAosgodbiqWuBoFjiWBsGj/2WnsyxtgqqMG+fyQBircht
x1lvo9JTgr/PgucPBuiEhBqwUbJIivjiBKkze7mYMSpPV9TkAWHhdd+KIE3gV0AwsaGuWROSIijH
eo9i08LgGB0jCDkhryRUvahyEFnidc6IkaMismP3Q5gDbpqV0DY3VvnyZQeqCx5uk1wJApfL/COf
dO54ePJOiGe7YoSVIp/9tQpaUtA/shAa2mRfBZAPQhLEA2hWeFHmASbujbrihKXNbtm2tk3onV1z
wLvH5/fJyyyCiihjPHNhPd1QCUymZSeFBGwekqXUPms5prUx2S/XZz1yHlJQ9KHJD8b2QzK1xeiE
AHMXoswWj9zowdWFgPFfW5v3OABzXG2O5i8zjAOx+uQ1d5pMYX+1FzYwCTq9crwQZWdeMsHR/Zr7
v8cThp3jazPySh7U7iRS3d5dDNgUNGCM7hGuVZgXueRTnC1oouKQE5CTHriC+TreKgJXAySLkp1a
h1trDKXdDeDU8c0FtyCmgUmKsPM1G9BHnH4ASTYD5cEQWmxs2AQ/1cHTp6Sih0sGhJLNy1IwL60V
nNgaURHMH2Hpydlm5u3AHb21jgvzeF9z1zVXoJ8RDaLsQKdFWyB13qbKo219qFSslYOTPjObdTgL
o/nMx82Ug74jOGV3ovqqPgO8bGKxpmx4QYo409DS3Cd3P/YRPREZfuxDGLn4WieevTO33xlImrOf
URqo793ZALkTxONbD3H+51GQp0ZNSHsZf59Evx68cqtBaBFjcqNkp/Y5nvGDcKZPb0/+htQij/6Z
wPQ8snsRewHzAAbH/nIa4Xn61loCghWpIS+DsfanISf4I98czYauFpPKa+cvU0tCL4DSP05Jjp4O
FsrXklq9IAYYKT+Za6L5NrhYAT5BP4vQmXSur8jZ08fUzsLgC5K8AqSk9knAKk/jEUDDr20VJkho
Wr7+m977vdEa/nxx2ftoBoN3MUPNeTUXwtjxLpbS79vLPDxx2kKTpw9UtzTuh98m6Fnvx5otkkeF
UOhV7JeMjo1OzmMXcjT5cF8+IbfuaKnoad3HLue4u5qnoLHN2ykJoGdrv7lGXYj4ytnQBVAtBZPx
GrK2jTm+WREUybenDi2X58IweQiBmL1wD5T0IROHQ/aKOtpb74XvP0sTO0n85siKXxJKjd2Y3P/4
bCErtXfhQ5O72c5oVRL4JwugX3WgjOeu8zHLPtGcQuaAb62GOtxzE/FXepXp+EjZOX2DXdXkUEX+
7X5/GKFZozE7uwYnly0OpdffBKPsT+eDIednTUnkO7llbethTfywYRFWFBf1BS4zYMviBGqMdl3s
FOQziqRcb1XrztCVYt0UQyNPfTkouE8M4WDV0pV8IUMtY4WmZz1kOK/8xeU1iNYYuPtUe0Jm+kCx
xA8kXYt1YtQ7EDQcuqDPofEgjtmw4VBYMbbPJHIC9xGtxF8zVrT1rTXU9CJIY8B3NeoB/ux6mQdA
vzmOCsPMwbW8FxSBuv/tXU0mmzWCVTztwlWtw21zMtQahlTxOe4wCG/7R9ZP/HUrwxAkCd+FvJa6
yk3urHtn6peOboho7p3+lFCPtl6iI0r0ei2OIC9LPwnpe7e2avAQGGFb9OT4XdrFBrUbsXxY4h6O
cDVMPW8kNPfXcV+vPMxRBOhv3mBEsGoAYO7TWN/oQ2nH9NL+8yucTvSNLWNMBsr6LJNItUbsGIR+
1tKArCsigHzGLCKktaE+hII0CqiVoKYzVc7djsI6gHfs6RWQ1Xuz7o9XMnc9ZvJskCRhv5PFwylx
8adajGUDOdxpT5lRlgmu+Y15zVx5ipTRb9MB/uM3xgxiKQDdbX4nWYl4iZ5Jj7O4UGyAbA8M91Gn
RGUcjE+k1/v1bAFLyP0ta0i7Qdtv4eZXsFXk4gb1DvYb8UHgInVEfyr02/H1304WP8uwSVj7hNr8
n26e7LXlWC61UQdp5pHY3tkP/MnkGTBdoB+xuEoPHCIz78nZrE/VjXSZhRBdE33pDg0699YbVPo6
xZekPntboT53aLhtfENpcpzodsD9pjRZV3Sa2t47ml40PDW8lOiAb8MAqd4c9X6Ksq3VMkJQFAO2
anDISjw5QXCGnArSB0/EpL0nCH0Pddhu9D/mKZP9B9X6BBKcbv65l4vsl822z4xaCCBpcMkSETVj
Bogon0UfrKVQSipD/JQAtD0jepKxf+NB0aqy877G+HCOvm8k4ZVUMO3yQJP+Bm04R4Tc/9TGtGNN
4rnj9SbrUPfb3cEYc72ReEc0LYe+R+Cc/isV1AyBGHgemxaeLKMC3UXsMbRuWhDTCJypOpjXHnu7
1BA9tKVcySzjZAOcwT6h8CECACH9mbZXHZXrfwc3O0+3JCnWUzbYH4ewkdEuASb0bHTMl2E8803t
tqvdNJKdNpUoBeN/dC8//N41qKtWTlDqGC4A3kr6PjqO82zpDVfk6Qu2uDKOIgFMAVYE5wmc6+Rw
HjY2SR+dvJrve/C3kIJiS7Pvk7B6gB70NCB2fj7fkqtmVEiS+6mqDmRm/4n+nEuSckp8IsQHF75Q
VPdlyGX8BAZHO+F3bpsI4T9hHjnyidBtC0r29KY83zlEqd1gSzvAb+uqyWFfRBdv1MVNMn3QHmqJ
Sj6t40w2sC/LluNX/Q/DVJECjLHpYJlqH7ylGZ8n0G9MLE8muwGvKi1nE2CWfR8BS45Nq24rMZCb
8X1e1jDLsBKP2VMa0eZYnGUt78ZrqrYozyfULhD1WNxp+g1UC0xROrkDjbbg+ctJTSIBBRnvob6T
MIzgC/1VQGURegETO4NryPabJbgVZao6cMxtsKPfxJPQqKo86RpoS0hrH4IMktajiu/mqigKb1xx
2r8Ux7Ge5t8NIpwcIldFsukgnkvydkRuJaxZXW0Un/tjn+crjZN4QG3kccpYSt2uglHFPeh3dQQ+
wTPo7CVhQOFETdjakZ5KJXrWlf2tnXlWFkNUNnJMHFH8jr4JY05Awn7h8eFzR30jx9OChY3YYRCQ
OZyoRLo/fDz4ex0K5sjcEREnwmT2hqW2B6kywbGdbKmIlykG3v/0q66blKEpp41NEHhQ7HRSnjmb
603suUZgkrsQQndafazCLHR83tCqNCLsFiwTowLxDmFfoHz9b24Rx1r8A5t7sePxQvj8mZCPHBqp
K4rbWiakGaNbKwlWMECYSzrAMhgkhikIdT8N54WDtUnZ8T9JZ+vQkx4WjAkctA8hMBe/NsC5hxBO
iEY/oiPZ4XBp+RNdKg3LMK8t7c/GVJbsVcyMU0aFV1UPT3zeHN9EFgLs+OWRF+P1fPbNDgiJPncb
qjdZlKW6SCIN8ddFxhE66t0U/wzoyVejvYilDk2UPuu8qWADTNs6F546zHzSvogj6mBhCog5L3iX
osRXrOpXYgRpkRUlDcsCKaWOmiR8kd8DM1Nh5oGm0iiDXfLOMIFtkQl4+OIXN2917zCLvs76JPoc
4b3rndqFTw5sQdDegPE5xKZiDqMxK6x2wYfECPIKn3mK9mKVrRADj1rdxEZXK5P/5j/vwmGT/pOe
QUMKHOnuW7j62/4XWTHPiAWe6vzECDbsMimYQGjhEzsnKB2FgTC/SLLPfIX/+7nfkELTxjiay3en
E9bdsqQZuccBIr4lLE/+STnwqK3LrK1LqfDSNC+Cqdp0ul3EA4T0Qqf4Unwc6lvszlicGoEPyOMo
YTW5odcCTowHc3XrJ1aWfVH70cMXjYMlDtnl+AgwoHv7R+ISA37XYz8E3vJ+7G/JhuD+gy6MNybv
zc4MEeNQftF+Jy514OtLIx08ewzsjSMYVDtXzoIG6irDITQ+OaME6m6fMb9LvMyYwiAOdwz5lrNg
MaGinNZyOfUSDv45pVqZfvc/hhIE5wJaFJTZKv03XmtpQi5DYNWNe4JY2ypR+av6GvQb6Sju8QVL
spo3JJch9droplsiADhh59MKSodZKumTAEtnDstUdrzPeHgEmyKfYlVoSUNYQ0PO+DmMYh2IRCqN
2uX9yektmXCdnk0pKDqOTWDqas+ff7XFUSOxoJ4bTFhbkeI11tL6UqhwPkISumOIocW0vyhW+jC1
WT0t1YQiUZ6WYxIDLHJcWvNqXWwPcPwZChOe4kaaqtgQEsh0r+u6cov6FENIc2/aOdx2wzp7VZIH
sG5Y9UYrYUCNDXe5ztEEhOGHT2rHjSY9mseix+v3Eitusr8LyxaryJ1iFmnDCELQ2IHIhsGTaqDQ
xtWDWl/DiH8yggYPg4LkvXWZz1MbybHVh8o31Ahk7B/B60eILjcwrVVCe7gJ0NfCv2S5TA6qaxm0
NCUgPAYxRgUFnZuascbQuM3U2/n1R9FYdYGtNib4mPlK9mv8DywKQDcv+KTs0jcPsvy6QbDYustC
q057D7aUm7Ce6KJUcSKaM3y1eqvQvsJQ5TL77Ohy47H/B7p79o/8ouRRRKP/QmcPKEmE57avhp98
+qixj2BWsC3dIhn/IW7G0dlBNhzFzVsQKnmmnZLQjLw0nywqznvU42j3jOk/oHM1qBZLJZ3PSD12
k1zi1s5gyEHNWgAnPq4ywDaqJ5mt4EroyZlsc76QlE84hMSeS5kahVBLxIXJyLN6AeHg85fSDda6
1ad6XDifdcOcl5Mx+Sk/bsrsaNodp9w9jyaI+8QWrEIAu3Zquhbat4BlwXjlp/EBcRPimxmeMe1Q
UYjMtvYUbqT0bFQqNg/LTlKhjb0YJxIaU2VItYNrzTPCxfzOtRF525+dUeiC6Bho1p0gkCpZ/iPK
NloYKAWytxoCrqTLaVJu6k+rNYhC6Dj5apfU7FYP3ScXWQPq2tK57OdhqvUCOa/3Xh0Mo8P5gYW9
QsvHTLsReCRJ7VUpRdayQZJAYz7JZYpwXU27fZUEEdoquQydFAjAA8DJtZUC0SWkws25nDafUN8G
hpFPVEUVvW9FN9KplHhfGU8AvRY8aVM0DAdLsfBMtAZhtHcKGS8UJPmtTIGN1kodU2C9imenee24
IfcyaPr8aRSs2yqF9fL9FOG2vzPXhCDDXo/XZQ4SFt1SBr5BeA0I/+4ERL3ivX9//1DrvendzoQ1
6ALHa4qY7ad5gWcU+abYu3nEA2mDcTCJK29pwn2Q0k1UK5zMmpbPWfsQRco8YoX6teFkjCxW/YVp
6FlfqnNykkP4NNUUsjQb44limcqZ9zKMshhqpvYWLw+vjhQBxUU5A78rVgkCItOpK92xe2dKplb+
Wmd1eA13gb2GM6oe4Gor303Tu1NjGhsOr23nTrFlWlnjY5IWC764oq/kEUqebWsFTU9acL1OgUTb
nWqdXl+SSvZ/hNM6p+53PrhcKBW6SnNhRbUqhjGeNdvWFms/tguXfT4wbibQmmOwCm06SoKK7fnD
ynDVgVHLIMsxSLWDt1NiOPUzmBHRJaVkoyBsqQ+SM2qjdKpUDJ+XUHzopBUs2lcoYamdyXkBMumj
z/2TveFvJxYdK1nJFA7VCMRnvXXi5e5nkNMquDbCitaL8SZswi9LR7jxIefDzkdVWz2Ae3Lr6RdK
zY8zAhWOlkL2q/+CZYN3/QcTx6l+pwXa9IRv9kn0YUcU+jGPE/zaTtHMUOzVO6W2dEezd9lFzKNb
YPQbmeDzT0lQ++Cf5Q7lfomyRdZR6wo0VxTrJe3v7MFrr5PlOmm8KRDDInsio3mAAmzVR34N4p8g
/k0kUvAHVGoney2cxsjIwCMa5TUwtHUGA4RpgP7zKs8eGtu6vucNdUd+egB/ZvmtRmaVCJYLbWGg
BHjkXOuFQQWsa2zArSd8tyaqzwOIj47pdPRlwlNwwt2j/oHapjddL4EeC35FDlEJBSuAZHVFVPQI
wV1nmIu8Ca2ZWieeWjUq7SUvvR5OYXveCrjOvKtnykm0BDxC9sQ/dA0riuu/6SaBksvPFv+w4OEq
jkqft2UifnJ35+VmUHMaGSRE15v0wpsEYZTMTc/aTRbRiegjqCFEN3kUOoTdq+mD5XRAOqClRY4h
Fu8e/pwo909vMXUBx2tJ9fI9p7hJPX3Fj/OdWhCON+Jeb9yKR9R5cNJ1tj0pXJU+gAF13S2uSRH3
Utbmrb3D2EyNO6q9MEgp+EvsIMBmbWDAPP2zItSMlQ4qcmoMFonMASJKNJJNzdu7VeRgpotpJng+
g+xXeuXrtaFOa/KR9SZVW+GDcnR5ir+2/RvuKVnjId1jYu9hgTnB6imjal/urPUrXKG1dbqitLO3
7fLZntSWC06YKyxLcHMHvYW7Vl5iJ6vzu6lqO0yxuzhpZC8kQ03mUhArPFwWEe2POpFpcV4kzlDe
d8ScEx4/KPoAvTYYRkpC+2Y4cJXd1y9ObkJwExZe+QPkGonOopSt+VoIZxgg7+FU5EvuYwlDTkDx
Sq35y7wJpjZ6ohOKO/o5xJEBpfYBvcokfdJIKj0yenxGWpsGLkVI+GjRogS9BlxSwIWYRJmJFuSK
qIWUw82qriuartJpFczovsmKctuD5PDli2l/LwWDb2TCiDueFtPY4tTLNF5riDPTMSD8wYgijJ29
L8qCXD1B8DbSZU16rMTMT4xQ/s4m8pq6AGTrEqgXRA9voqN3kTatFMMRjDNni35rn1Rwxr4d/jC/
NUXnvjGulAJ1WVTmXrRu4FtdffNu6+pRfax1I/6w9wsPxJ4JvLHiKRLxvbi8Lt2Q3waTK1inT/bi
wmrQqvmoMw9mnE9/p/7Or3qLfHpe8ITIwn4ItFf4SSZz+5AJGFXbTfnTQhHCcqEEQ1BI7l86mRfs
9WLLW3GpcnejfkvnYytIq5F0g8KVwu6yJahGy6takj7+/BOWe6TOlPYdmJTouQEzmPMYRs8E9DAW
U+U+DjfmLBKFD73pjGGgnxVJ9IJWIT5wUTlLm6ycLJm56Pr50yfqFm18qJqcrb6QAlvg6i+exU8Q
7POg5ZiEE4+TDEFX3OwohztI0yIXz5HqugsESTXy+xOd/bfK0lKH577xIipF4oy641KycUkFLtuC
c27R7RU6CDt/kLfyrDZ+763jNoB99lxeLfGTY0sVl9SHz/nMnFQBv2cPT7UIAHC91t/afsWsiBK3
lLE9cepr4sWy3KuLgj+sGuAmCXqPM/khgDxg8Hki5pyK2wRjETD6ktpLDqRGWQrNEjRAy0VAgFY8
ruQ0LccSZq0KPpYQe2Nokhs9T3nZSkPiAyNJYQJoPTVWkNR7hUWIUJVqEjbiEkvLxRQ7wEds8/1e
5IpvbPSVcC3Lk9LSGGq7v2DzRjZAoZVgroJ9oA0GngIC4TKXXespMvzeMo5AJR8qBWGoUazuPc5J
13gbhbz1y5uUF31vvzRX5zOttXB4RKuBryVlKqGXMOa5DT5FQzQdho7PtUBx9GgOxZnxk1LuM6gS
2nlXpQDmOiPwXUXqIT8hkUR3rHHrlFl4bRkgl87h3VSjIy/u+NKxRknVxEUthUVos6FalRZLp0lI
yHEglSUuZ5XhnpwWX8cUkiFx92EGA2J8h7KfX+FGxkvvYT1eNDRhpoG+FMWX2HTFHFN2MRgIxDBa
K1sMDnB+nqYTRspfj2WPVMD39B7Z4tEwsXFkhoTlXtK4laa0sKxQ368/e/mz/xbK+41GbWznryDF
2wZ0W/fLmX+75AiZd+FwoK7mdlOQ7VJsY+jPPoOTG9RGp1oLYW1rxaXaI3rnme9tGqFfO5Rjt6Pd
HUXA1uFk1dIrq33RoSGGWo72wtk7YIH1JS1hsK0H3q2dkaS2CWg+B7CxYnvGQ2z1PJXHUBrLUqKB
68UITgrXtOw4+oLQbCFi5ZausoASYxvBIGHTjhQk3g3V6w6oYGP0pEt3pCugBW+Rze2vi0bSchD+
HTePuiUmGK3JgurfJvWwoCc1iBFLGMe36UZs6j/vDR9qPeeTHdF/HrSzdWR5YzXUqhHR5SmwyBef
xd6k1/EJjAugJ9iNjq/HGIai7eXo6z+x+saTFBEQXnmy9nMF88rfvhr7AW/UFQ41EsRqOj76JmC9
WHfWyFozvctvl+sZ+X+yaS7Hhxuc2awtHdDaDUF+D8CEIiuSyr8NkmQKQbtD7G040Ux0avLXfJ2w
slJTZ+q/EYyTF+2A/il8KzuZVQyiCqgTCtOjV5B+5Ku7e85CE/FBt9mIIiK9BvQaoAM8xgU7a8jX
KH9lRdjgk2tgHlr5yE7C5c9mNA77iE+D/5UEYEx6Cq2HtSYlQB5MuFnwPoNhS8siCQ10VZWR395D
c9q7HuiKgt1hecS/I4cMcbr4BRF/n6deiyMKZckYu4aei7KFixqnVWa1rsG78AfGl8Q6p9CaF7EY
zBApEErALR9GyFQY9H5ZbZRwH0s+a3i3lNl0KGdoe+fEgNyPUM707EuCkozwvyJJkZ7oFGZh3q+E
kXUHdSROCcLVK9dcLW8gzov2KG+gPEVnA5KfOiuqICGtizzzGz58Kp2gPi6L9ECk9j7afD1B73Fe
NOVgRp2PoAbtEUomR4SVYw3BJMNSmYuy1LU6DVYNdF5/czSc9ebPbbHDcX+XVOiVB02BMNiGTwQR
hXfBTwhMkdvByliFW4wys8Bmw3Oli8GYZyMiUgzmfdkQ7jRLah7Z9ZRl2gRlGqfHyamR2h5Wpsa9
wysHbDbzYtUg7yeoQRQGc2zYGSqYfEH+AqdsbURfprGltACJZYvw03vc/xCx/0Iijy9ct+to2HLr
APBnY/eg5589GEAxuybtjgBWeGF9Uno9EDo54JehR5/Ow8bWYmkI4wVryKV8s/5z6oYz7QJ3nTQj
qdVJgzcNMu4lN9Tj61ueGyBd1x3mNTl32SxMSuDT1zv868OCqOTc22Xc0hMMVdtuyV/JeEnpeHsa
Xc6Byjymko8QpTJthr8KPibEa25Ya63Mx8xiJebShtZtUE01Rp9durkYYE8Yig7m7pQ/u9VSKOcR
x7N+WhxTM9tM18HQ1TUtaR7X9S4GxY3rnIdvl+EOvq2HwuvM34s8EZ5KUYfR3KHsWPQpxQ2Q+4Gq
fJ/Nk77hxuZLhceXOz5VFV/7i+6q9o8ZJrwPjSRR3BZ4gdVdgIOqiPl/9yD3F6MSoYU5DkRbfL/l
lelKWYT4NqJSuJ2DSn5tkFLsgvqFZB5d2Fz1ldAOuqKR/4GlwgeyGnEzbfPDTY0AJC6tHdJ9UBX+
xOlef0dqsWgxPWs/LgKYodb25Xpe9FSt5UPAgQ8lkGOZBGBL1/5ot+/RBIjOgxDUcFQtDhpbE3+U
SgnAZAb+nGpfjdCQmo4v2r6WKC6nE/DQhYx+Smyskx/y0fytCgi/5fEQwbHnHSMCmUNI3/aBU/e/
4+sfbIlkoNBBvFe+Vl8C/sqar4vkVc4F8ITmIg/guAkpAxy0y0YpTL7HXAilsHjDHI+FOC/0Ab8l
dbRSvgGFi/tnD8AMthWvSqhLslWXZyHzQdkWEwhr73pULEnHwRVpnYZmasG+xV88pyd9dZCp4rCq
54LNkSzEVo5gaaFJZuQIw/RkUWMdEjpHr6tGIyT4fW/BiAmcXaFREYdayv3kxg6YQZptabbyiAq7
DEEtQEQ2wFivqY2fAq++PG4nkfe2w89LR2fu/WSJOpSLZnHBRQlY5FdRE/wpyjtcW3I/PecMHLOL
8q+MXlo3yOdVgfmj4yXjVvOAsw4hJMFZvY0z7asklhhmEGIDmwIpuydagpXdNV/AB0ZKDUlrMv41
y/YjQmm16roZ+fJanQ7rx3NFQMx5EMsdcMCyqQdUi099pJB7Le/Jx2NDg4U/rMah9WlmYN60/Akt
oyahms10h+XfSgFS80PapeaQjShoVI99P/2aaAar8l3IKB+M3qluHHny9ATB7KgL1twhweRTObCR
LrnnaUviWq65SLBcPNVavkrvpFqrCgiizWOZJux8aaqXkh/CdWSL52Flbd3cRPyhh5pRZQxAyYSL
mDj4ax7dBGOLDBvjO4LFwmc4bSqK5l4Nt5Wx2zminPCsCYEzWkgddxIonLld/ZwFQ4kfw9/XtxUX
aWzmdhSusKuFR5kKJdMHRIViRN1chRnYS0rRpddy+XlGgKCJneGFbpCNlJ1FSjUjqiFCHkTkPf+6
aOdXTgofjt4ldWR7lZ5l++8qL10/PBSzUyNKvPxNi47WpSKNjOODVhuju+cmf/BrQonFaQqcwVCH
bBZRJT6woT7vjRE7a68Q1iKGZj7QvddwZctQladO/50KfUMGme2DltI9Rp0fAsiBBL+8NKs8YAfW
iJ1Hph3XTckDzfaI1irJJtpj1uSoL2NSEFwzSOgeP8dDSg+L2Vtfl67PebOfyd16T/ORrdePVQYj
1TxwA0LR47ac5lInQSU+7JGI9+DBbjJcw6yn8P/xYNHkGk+DbzZG0W/73FRGwcrSrfydQu2wjuv0
YqojeGXh7VRMyHgVZH00lqiVRo/Ok14GSu8iT3sqSdC0hpyFoAmVRxS4kpDvEKq6+JlPCDrx3V+p
KMkPTk4uLNvpa1xD1gcyYeM+xpA++WQXpT7GBolfwCUXFuR6FQQIP1Od6SAV11vOplVj0s099gC0
usr8dqKhWqQvcLpLfgKvfXuFGuZLBO/rArcwDym4r43fGhFHVmyv5lfsZC6UL8mCcdDRBvTcR0KD
rr7WFUAvKRSsrdlJm6pB2tbaqCS0BMOgeH9n6PEfMpNDGVPH3sgs/Ya5G0txnJ6V35c+ke3Sk752
Dulq1WMD9xoa0ytOBy1z4orgYuEoVTkMMr9W3yARVAFQ+jDCFLEAcSf9ItXZKddxb2g9f0DhJcs1
EZ+1a4q2CNnvMgdWpvKLX7M+KTscasqqvob8lcbgLXA0akoBB6JPOuxLBAEp6eMiENfXEEu/HQlr
1maahPhtcJWlnL9QJDDUX9giYnAO/05yWib0W124tIgtNLttXJ5/nSnQbSjxT9qU6ebKuIBAVim9
qYRc52YK8+/CbwcggslA/StTFPZ4SWVCWvwqVfaZSHUOLjl7YUiDVOE/OAtBivaJHUp6kqkZuDo8
OPqq9MoR4+Y2SIhq+r0ZDDIqFZdWlh9p0V1M8ja8f1rGNc4OwJdXrmDT6H964P+mZxoIkujDzmQS
dKl80AbZ0lpFdi/3Stf2Yr7gTsWescDyT60bICEVomhnJ4y4Vmykb5sgv6bp7H+so1eP4e4192bx
OLtO5B6zFSIzWRN5P6yvdn2gXNa731KkguTrLvI90W3QlvTBj/ibE3oYbk6xIhl4ZLa3WdHfG8/d
HXtHk3GLrpZV+9vxs7sWc1s8zRcvxMr7J5UkZYgBhUp9ROpDXBRIHRDNU9DnsegFoYpniRLTlxfw
2mfNLeOih4B+EMnFmvdbSgI8sW8gyFlMkv4ygNOjbH0WZUCv1SiMiTxgkzPaNE1PqsCcIwoeGoT8
9YvS4eRTl+DHQvOh99iCyFC0tHl6EHE58KES1WRDorEy05ge+XtW5IBqcrOi6wjnN3J8F9iHkZWQ
98FjI+B1T10YdaUX1yF1JZBaEBZqRCFiSHrMjpR1qDZ1bFqqx5mDBMXDx+STK+oQRNid2fF54wOB
LAlTvwmoXT+IlnGWGl1oqWMPbUAwOXW/+EYUIQjGmx9FI7udt9QHu9sIc9lwFs8wxkVW1rPCYy3c
1YIkf4QPFxAWK/JpSJIiNampyQ7dw0p5UlcSCnvvJuKxy2KWWEW2rWMJKDhTHwfzS7gN3S2li1rl
PIs+M5Hq6v7VCfU5aGQ2uxGx7GsULB+/A3nZpGbrapl43oROXPDKUEgZEZ86GUkr+uQ5g10uOgoz
jBOklQAMeRpTkKytppD3M/tO7XVDAlznUJ59TqLKJGbfHqOfteYVXG9qKzabEqp/mS2B2+xSylkb
lJ3nhS69iSW/syaMaruisxXwQrIPrVxxsOAwn5h6pSfpNLkoA6gFoe4J94g0DcQ12opTef+iKlAU
Qmc2nKSFFd1pWDHyo+LBwfM3TrKSpJkizMdc6TpchOkskw55dB/4uzFkDkDhTbZGrlv9VejERK2r
t+HKju8S9SipU15mgqPEm8c+FvSCy7gaUAPyeDsDj+aekB+dEMRy43qbi7d04FmsbQkOEQBn7EHA
P9aV8Yr/D06DoXR8Jb0AnyZ32uAKJEh4NLdnHX0g9ZlQMsp1jh1abyfEkBdQa0NhOi2yzkoZMdj1
pCM8Zfe3jtUvinmlKBvU5JExYXCwXrUoYDXgUpexKBDR8Na0HCJVRTCHnQXsqphcNPF+8SHn6Loi
G1D8+Mmqo1BSgEbIwU6Ozet2CrZXBMLyIaNzZnPWOCkDr70Kmi3BX4il3wye8Qmterf0n7Nqp6nY
X4pvQOKro/+C+FFK9n1bD9TZ2kwhnzcBHBfKwrFqZeurFmVc34A672VNHXh9sYuZMnSI9ehpTfZi
Db/+1LPEk39j1Gm7AnSLTWoTHrW4Z5zZKlCbOzLBjH72Np/Bk0j3lpjt8p8nQnw+b1pcjcrsi7dz
aJfaG18jbGJBQuUEgzZTn2lE+NXqB6pF8SVtO0IZZcFWqzHDjhaSOJXdV7ZeI99l7sj6Z2vlJO7+
d+NqNUtEzqWbmyzEt+pv1de7Zh+JehlEmlHM/Js6YQ9ms0jfHgHuUuqi4Xc+IdDB3XeAQ2MDPjyh
KyS0CjSVN0tf1p/7WYeKyl5KRsGegynpoBH2aBNSeboZ5qJFc7grsr39+lF7TmcLi4Q6GUT4kwmx
80YnhCB3ioRacgObyNL/5iQN5SFU3slonQIL80FVfCiCUpGO+KZDiiSpUcFFyTTBqdOzdcJ4mOM+
i4E8709SQvnbmsnmglh8pJKmEWeb1Xe/3sI656UGQIXytPV/Kh5eTIn3RY0zSpFhv34nRArKo9b1
paw7FsQH+HbKYgsOr4TXDDCEeaw4q6Ovo4TdQvtyEA+AdD3ugINB2ZzV0qJi9cIsaAO2/waKVx+S
GUj3sS2xru+iMt8hzRRpcoVwysZ++s7kRvQ4Cc1SXGOHYW6/Vb+fS6aPnJMrtaKppextnq0/zAAX
wLbbotF/3lnNfkcFqA1w+kh09pfP0GdXtGe5A1OcwzGAtqCD3CNJwr0kFaHgRrZ8+nFg8WaWyQ5c
dYDiStVwYPhZqTvXHlQfvC7SnuBlmL9Fj/mbXMarl5tzi/QNlny12VkFconBmi/hnz7s8Xxfltte
zHheP/l0hS2kJOM63h0WdZVLmqcYf49Ba7K9Em2pZaTinKiCJ/cr20ZYj0OBVWk8PnqiYOgqJN9D
21JefBpTqqjrXiWiB/DtMn0tZmMQ1m4Iwc3FERcrr66ynJFyttxGzTnRisWyLryOQdh2kYnemTNg
+jUFyuC1WwG5OvyQBL0qwpkvXGiedoBpgXi6BBJKV+XQqEE+9uL5Z63BQl7tMfwKJl/LJ3yzgUTj
Re2N7I3v5AJG5LIQCfP/beguY7xf+jtqy1Etb0hyxZ7H9H+kozzJDkNzIDz1sbmZDH/cUOsU+aar
ZoNZJziKqAcDbBV/TUXMXa7VykL9oxp/xl5xlYOd6W4IGYEnXA3tLIfv6LdEt6o2t5b0O2h79LYA
zQiTtBJP4qT8zSU9Q2MMNiBlxsrPDnbeagvMul3V8HEKhezcsGon+0dA1izv7M7c0O7n/l2cnyc+
4LOqXkcpoyi5RQCJkn7gJZzyb22VqnE4Xni4yx0H/MwAmhHzBnrzdhF7
`pragma protect end_protected
