library ieee;
use ieee.std_logic_1164.all;

package root_package is

constant c_refi : integer := 10;
constant c_rfc : integer := 1;
constant noc_latency : integer := 2;
end root_package;
