// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
1g2rnxiFCNI+MVcCZ+VNFMwlI+LbkzmzmpH1XVo5AZEsdJm09MFjT+IZdilBf4M2
ewmkkyobgDICH3aMbjAlQ4G2xcOAg9nsPHSlATW0SB9+N1qMam/wepVfJdzlVLi0
V4eB6DvS/iWp3TbGrE8ScuHbn35yTn+o970mP4ZCNC1beI986irGmw==
//pragma protect end_key_block
//pragma protect digest_block
Pvc6M7xkTA/l30MpB3rE77E/AYA=
//pragma protect end_digest_block
//pragma protect data_block
ZD+GcidI8WCdmls31aTxNtRMkDOAIDTggQ1YptzVOMriC6Av727LnZpOoTkgk7k3
/kk5viX0hqz58Z2r7yJOOpiUDKoOJHPqg2WX1iSocH4M+sgxSkeKOZzjU61E6vLq
pc3HSVmRrZ6D0tA7aoHze1fzIetN7w374etHTB+bmMjZjevZxuExYTrHkbLUhP6F
k8pFVR2mHC3nsQ5lMMEW27CJJaMqHtv3/fDHHA8AScpmOg+BPTXkWBhIspExw65W
iyoob1heYpcR0mFJYNwG9s8/0EYUMRktGn8wPAvK4GXiQUa0zBV113lv5Zf4DGRN
RKssyooVhAdGJOhuFopTAPVehQ9+Gm72WiehIFJ2+Xr+FOhiizk1ZB82EzIASE8z
ZunODfhPD2OxY1HP3hUnKMCn8cIpCHkJZRGwOHLodGB7JifY9N8+tDL5TEida/eQ
4VXOK+SaAmvTGBktx1Mvzxw61a4OwkFCCH5JApnpV5E8kYsf/z4Ho3zWhJgndMDn
6dBzhgfjiitZRgwptaF03eknGrFvoeK0Sh8B09el2ulRd08Mg6pDvz1FyCLLzie7
zc+OSs0ddBAU23djGEUGXGApfKiOtlV4BmJi+k0NO7A87BqmJ7kE8NleHSeNR4JE
AA1j965DTuspxiF3E5jIkMfIMxZdHgCaxDpAf1PulYsfRfUJCCVKCNkJhJRQSAYV
lfg31TtSfhtCpSxCCfKFaTAzFmAsGCFKV5HdZtg4GYpHc6K6QfM28mruu2lgr0QJ
SU51j79+Vj1ebl9G0wdrjlpp2or7qb5z35uACtW/SI1wTn/JYI5C2KX9XutWO857
2pqWf2QQYtJN+TLjPKULWQ/iW8U71tzvhAWniBiimJyrTwtMcbg84D99bwP/W4lz
M7SHZ4rFdUY5zXPB+TqJlPs6yaUEL77ZNyHPI/geZC4ka223SNNuMP0FyyaTwrEs
OKPM8E2fndQisBcw9CQ8minypeBrzATfAEuoFbQYbrcYr3krd+d0oAQqT3w4v3JA
cAxtEuGuQnPUth6zUJbIafN/dGGrbN9EZ0qScpiE19jFwabIBsvO+DyCqAhLMCsX
B7L3zmdMz5MT+OGbCTE3VgULHmSIeCNzUXqsY3BFaYBmDiYoydfcojm/0P5MXzN+
DkOWC/+945xHfxD5B/gwpNwh7ruD1TldsmmSn48aYEyZdT89AKFr0PbB5P5C5Dwb
Fl9ARPY413GWijaDZUTluE0bXbcrJvjTl/etQRqjE09ycqHmq3G98KiUxeDqA02l
CUQmpQd0mw6MHL4drflzmUpRp32AfVfUPkxwVyOQfHziXlS+S/dA2WEOaRtpWZZK
nyuc60t6csU8qVQJyA1pISIyOxQdLlhiPXl0HssR+x6m56jfj6GDJmeTZHHfrqB3
J3/r1YjuLXZ+xwsYyXnQy54s895KmsoAr5Q0mor2oBE/BjvpPtXcxy+U2QM8jYZU
5lo/jBZnFENZHTUCnixxbVNZnMGB3e+tBbMKTpquqLfmoMUFxAhlh5LLv+lcKkGU
MpZ2g0EI3lgJZm+9Mbi4ELLIsZYwFEsg/D5MzHOISPZXJCsC17N/gpr+lX0qWF6P
QHkhXYg+vZApCGCegQo+dtbQ2ZIU1JvPxf5BzUsx4rHSfaEy20DW+DvOL/hRbqM/
mNC30w6+4vCFkzG2h7i/dlk/wEBza47KLTTEQt9TrlDrkSe/ZQqR8IoBh3B2LCyY
+nL3kw7IXrQ8dp/AoUAmFKZ4+GtpspQXndhTafaB4geE9hFSOQkmDk99AjPnaw4K
qu3x1KUrqn/TWXKDWvKP91QtkwGQdU+YCkXc/V05llvhvjkEp59wzsnz01qlaXZF
GW2Yp9jq7vVM6eGUn9MR5e+yY3Ga4YFjnx20dv8ObqzJ4x8z8HvIARlROvHwdW9e
c6vj0206iC4RgF7S4ORgsuKauF2NvbQIwFklsRl88Wr0+CGK4HyTwHroHZza9/jv
h/kjz2m0vsY2k/a1CN0dFyynUjXyk54GamavBSgdjCMabnWf5dQx9fESkvzQZupm
XhtWAT0fLfsCJKCWcPBXmBHWxL9H2vWlGZPPapdo9/hTL97wHjR7knHzoXemySx7
ukanaJQVE7UUU0Ng45FwUNmxkILL2a2u4ccTJEKr5IMcg6ajy05xpojV8APEmtnC
MG5/cSLPHQ/3dS9mtbPOTyqXJyFPswa/M8e7VPvUG4ka1ZZka8aHNZSn2fQlsn6H
jYlaraEy4g7DaAB91Mvbw4tI5/NXPg4J6N6WZBPFGZKEnrhMAtm1+b45qDRTRv6G
94+PdHjIZ8Dt2Uf5Jv39vCTp1xtmmoS/jg6Mx5N6fXj9upNrg+bz1Paa3tAPhmKX
oM3k1pHkwyfeFLeEnhyt4tyqGc/dVIqnvt9ZHEtZGG3lo3h/uhGkntIqsP7RUPgv
M+xQdsObIgsx1dSIfJxPraeE9fzZypP6SayJOogTySXZxGxg9YhfcxqVnH+WCpAW
xUCT26W+75VwjDzOekuTOoAxJPG84ObwYy9pJYJyGu0mTcs0qgrzlb6QlUNaGitB
ZaHSWHt03TJgJQIelgjU9oG3F5fSkZzJ7VMzYCiLivn0+tsfEdLBtYvDd3DjjrY+
VLCwLRnwEHLxR4IHrvhPRO+TW7MKKOGNDGnI7kTKx4415l5y+vEclDzrnRBc9P6r
gwQs+76PM1u3f0RP6CHzWmabkxIgFilYsMGHa2ImSRDnxqi1JMtS+JJeHQ0RyQ1C
SYrg0WKI/VZsMejQAHyM2eNU0n37WOHMuFjB9OVL+m9mkHAp7rf2L48o6nt6sTFc
k7xAqASOklrzO5DUdhnPiry0JpMiccZKF4xfJvD25W7GBms7byWLKBZ0vaKuFr0w
J9GakdRVmwqnQabLup/RfIc6D0X6C71CP3SOGj1+rxLIbi9CsAK+SbkUjpaC+usR
9y1fO9turnMAgBYlkjyfW6UL3kcOP3Ek+kZi8ZIh765HhOnY1T5X+Y8BVcjlbvdg
2JOfZGjANe/lRW1bAn3VOtCje18padNiuIE+SRELPGZOD9gAiEE4gMfpp2jlrjqd
fA3RV3Io0PG2EulXVp0pabm8Nt/m8y2ZxXz9zXfa7aYInEuZI2vAtJkKQMKnV1O+
MuVN6qQrsX71mhZFarSejBlTh5yNTyU477unav9quhcMQGKzGHELTx7mK+O47a7L
PNrag/qPTo307FtDKwEgmwNrfsERiPFSIrA8I17GMlRf/XAxCjCs9fye2W+GJ86G
mtKMS3grHeFPJXIjHvSYcRYOo/OYhBIigoe+kDzRMx6suxxkfn64BZWSn9HY36or
6DRW8ObHxyg5WkUvM20vvXiPD1o04VshwJgTAdjAgkBFmlNmuZ18a23bdF7Vmkcu
WMprZVRFKmk7Z2XpXjvQrkPApL+zZECSVy1PwXm5hhGle8Wevo9bwso7qV8rWyC7
URkVQYYIgESXdJGy3sqkJIi6OIRdugtr1J6EasKk2RCqeBw15lRcvtxiZL3PraNE
QDHh4e4H44D2wzqxZUNgKrEDnOrMtYL8hZlbuTh6TThhrl8/mmbJ3K/M80/Td3qd
L1qTVeCaNi+i4cebtT2K/8GJgMipksGrTUaI/4gAkkSGXREqHhwQe960bM6UYohS
Ey7Y2EKNG7/JZP22u3e/Vvv/zHHAsWZIrJApFdvThvt1WrlV40JeYxYV4IwmUyRy
6G/Rq3Ttz6xy/eQCkMrtZd1AxexOXDpmVELbU4Uo0K3Y80HZ5pLeVilD0XSx+lPg
sxoS9g8RAFcldXrTubwSYC6XjRP+PKHOWHpW82DAY1wG2hga6Z73Nu6TmKj5lWqi
nXapsKzhdVZW6eTPWc4jsxCZsCFw+/YrS0PJj1Tu1MJFZiNhU5zbeWzS1dlLRk0v
aHcuD2I2E5QhsztNNpb17AISYBrsCKussfTtH35e/AKpQLBg3n+jlWyUroFOFaqN
pDE806I2hPjN/h/NpKuF4Vw47w0vmhKofAt/fUaeH3+fS0V14IvWIRKijr8Yy2GE
efLCdigS0fEkdxT2MwOZeEVSHlaZrW9ga0JSa0FkzOUqy8UTsJ7nQsfSngR/i4HV
QfPqstYP1NH1YRxEjpgqbo9qJxJZ6NXxMQarz/e4sBM2ToOaSZ/B4fxXDrQxl2hR
31b2S6h42GUT0PN+F2t396L+Mz/Q3GPRxNH3RQHl1qGeg+Lqv+BVZ5ABvAZsaIMl
iX/CX9IyQrWvLXjcUkWrFCZqnvakqCYBlj3NHpxdUHWvqRrT6BDKyvuTTGFsq7Dw
2PcBT4xPweEI5n0q5c9n37a3wbYws2216HcWiDT5ux2LyvWpEizH+d7zZi7R/Leu
eAnqzJD7gqM9RjVyfq8NFNGrGmFO9xT34FGAT63Oyfak/MmuXfBm+152mItdbwuV
L3lXFp92FwDt8F8Cp4VBw6XnPKBb/Yxw0fELjlytJIbGvwN4Lg6zLnpC/DNW3seV
+Lq9Eh7J2JSHohVq/MAxkQL+t9VPI3SThuDTHsYFEZCODD85HojYvNhS7PYDXXGU
AT4YEWTsL2bjd0aa6dCmfNCXqRaYSyKFrOD+MynSbcPc4+YllblThf6DGuODwT0t
iv+6qj8/+vRq33lNigGZ/SRNbaLI/2ffFCSz/ceThRU1oGX+zzYk+/nR9zbo8zwk
tWKQ0wEoE4zIAbZxe0IrxpI0Ue0xGgCGJ0ROUinPBXmASByWtKg9NmK3PY3pBfv/
uuqCjFKf55dcIDMcBnA2E1In4t8oLM/akk/cydt4JXQJFIY/xUv/+HziwjQ+Az5Z
vPt89+LBRLrbSPxOdjKB4UgEl4Du62G8evIaNTpJi+YKeRPaQfxFHjIQYaMJNmRo
1gS7HN2SOx8NtXS8wATylNV4GI1vgkc89pf4bMDkdUDQGo56NtOKEgjBbeISSYrh
kb4YuEQaHjh7SlJy3BrZ2JPQCxShcaF5aF1+9qiqw38dz3rFnGjUIoUIS6bZM5fU
7IXniTmBsZt4d6v0qdDCX26mJkXyJFNxH+4zlS7hFBHq8vmERVqkrpwQNmUjlGF3
/YDNupLNpdNzhc0xDpPBBnG7nZyXaUHV6MHNCeLAgC1W2xwL0mv9Ik7nWugoq75Y
QPL7r9Ahlm5+cRJhyflBLf61JsiLK1GrxyH8fAXre43pI18zT9I9T9Ejhj1lZHl3
fsNEoi3QT9GqbSBaa+9QJzMFVff+YicG5CqJOrLzl1F6xIMsCIDlnBaFpSaBjuvG
6/2fAWvOUJIuV8nHLaJ3dyIIRXdvQ13VxsQm6b/AjpiYJSG/lUDHKz0p2R7VhSmo
6piqYrZvYDEw3TCJz755dt/zojxj7Q4jzABelFONMUqu9Fs+TEZson/VnRZB0MUJ
IuqXQB4T/LTsBrma/xPNjKjFGypfo4Yeo5T/XZF07fOKTVG+YR0eENgp+w/LCeJ8
1+JZUGbPRMaOoajweMeZVM1ZpS0NdQcCJYNxoUXaSjvcEg+OZZhx7qqX42swI7/L
L/o8/P5WmwS25K1dD6QhEJ2JC0ii0gnxpxsi5lkYQr5hu42ANT4+ETIdha58n4Om
zj4oVlCKE92FpJ3SEBLZ7EQLE/UXSWeHifDfxv0AjTqpSodX/rzZeyZuVWiNUdOJ
JK2T9qtvvjU94jNQU75IQbCf/hgPoxuLIFkYt8kSzDcQgQHKvX4LoU/VZ8/iGlUO
hbEiucm1AwynGOTQtdHMpW5QOGut3qTsM5dS3tHtWN3XqI0Icbo6r/XnO5UbKedi
nqI4AkOWEbjaWNTAupEHp6NM+3hxdYj5mntvqPhcuW7y3KlfGM/2TF4dZDK2t8l6
M+3SKSoD1mivxEZYMzKPviq1HwBZIQm5fcHSBH6HJdX3Yi/TbN4647pALz+9wAUZ
Ymib0Wm0GEMFLWpOtJswcFdW8GxE/ijL4cQv+eE7+OM5RwEeS0WEE0/7c7uX1Aeb
BvrQFq91wr+O0Y6u6D9tNsYvuF4aCuqLExdy1frkzfBgeOC6QkJ3/uMtDGFZP4HW
VKluDtJnirghSh+SzW4gRcYeZcosHADaLS/lFAv6tNbvUUFA1agYk3LN7Cz/X8Hf
QQDrcKs1ZrETrJ+miH6uw0oe8GhUhtUq2LE38LYDym8d4HjRzskc2NayP3CJUQvL
1TCMGWZxXyZYY3uJGlmS4MWHjWnlrZt7JqiSAVoAl5T8ewE/X95LPu3frNh3AK2J
WgS6Tljm152wNm11cSg1phBTxCuu7MotpcHEVLRk2vYCxAAtKVuRlYdokAu1PrAt
I+ZFHABXWepDCnkyAWwoXXixowsCn6HMti08FKYTkDjfh6vyYEw5pKZp2tVGCKY2
d/OfZB4AKU5ru+MfiHHc/Z22k+U6/lXICJ9+FfNBv2pv+tQ9weTtbCv+ig7aPrBc
+6JSgbsZBTMEsLTLSb2fB3NwW5vr7oSM0XQ9SMJbAyz4/9IxPtlnGKoeeAMoxIB1
BaH+8b3C5STx9s9p19BB4wCPSKVTEg5ranORcDgzoccAce/er4q0UkWb37oujV4Q
ISWsoz9XaIl9KAl2lGEqfCj9wS10UzOdcWYVSbmX7u7o/Yo8LaW8J6hehoYr7coG
W0ShKpKhLLbFJOde379j68cFLKpVek9Jzar0+Q+ztNuliXHkee94r84Yg2wzzRmN
G5vQR66SjhPwE7VOkqXrM2qHxwxvIXERCqbKDs2P7Tl11qMHVByD+QzAjMgcFbt/
F4uT0/n/mNIi4ECWJWIIREIlaTEIGODLV/oVV+jJ/U3vEvLxP8cXVNRMoFuasDWu
E18bkuguINhRvh+FgwDJ8qtlD18UmtGncEbRji11GG9iUKqmDGmL9jSiNL3jPbdW
0T+mM0GvrY38zZSTRr9wukCGd1A9WCAMyLQKKXfXqzV/tXh8Aev5H6Ioq0Q/8dyl
u9YyiXE6DYvf4AXbcZs00azjIT3doW1l1F16My2s++7XhpKtefujIBifJfn6wTUn
Y2oTqOk9tKFe+wcPvINbDGkIwZQCxmalVbYJaqWezJOuqFHxvJj7J1nuJM+CCRyF
m3Rg2BKrFD3dJWDReBgoEtqJTIZ9Sad5NlZ1CqiHwc+Zv5C9StxHlUJjX6YTYolC
VVlQno6fuzKk8n4xtq1LwPQ1HcN23yoq1aGUou+ZqBICO9nb4MDPCC+HNMSbU3gs
czK3rDLZCSE7s506yqkE4l/Yr2teWISlVlql66mw2mgvx7a7tyPUOMJKQRfww1E1
CjOQWbvnii8LROwB0Xc68/iD0VyaGXy5iQtAFkq6k+C/zK0xCg0pfBhdr2RSjkAN
Wz9gJ5tI54eU9A1BzS/BXnWefC5yGavtVHgbo1GGkOvVPNq47lv7ho9bwBn6VXZ8
85FZZmdmJTOxF5dqkwVjR0U35zx36CdctMwkdgxu8mo=
//pragma protect end_data_block
//pragma protect digest_block
7cXDTFHWQ2HNfTKCCDGz3b3bL6Y=
//pragma protect end_digest_block
//pragma protect end_protected
