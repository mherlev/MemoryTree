// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
q+EjAmHqUmow5oE6B4PZ+5N0lyQc3DlWtgngOY7AiRFIrCWloHtqGUB5L4KVoGsd
2LMRqEaiqCtHP5kAGws23FFM7/QOpgYezPhkreOiCVbA9NOfVT3HP5XYq0q1I1fi
ydvd1qBRagiZUzEUmxwl4DfjCAMm5cG28CXN65VTCGGx3IkOnoYJHg==
//pragma protect end_key_block
//pragma protect digest_block
0ebIAN8VGvGMDjwvIeumzQyDpak=
//pragma protect end_digest_block
//pragma protect data_block
kDbaUJPMXMOHqM9jaoNMB/KEriAVXm0qeeW0LgiQzGxGqVPhrdxnF0VyzpBpWqbQ
UvPV3nMfHYodCedsylotramQA5wsh6oRTuWaYHiEUQTPj799vmD4xOhm0HyPuk0m
bQIhgo+Dv2vgbi6TCsDyhvzC55vourzqF4oTZ3QUHn9N6FASZyJoj1udwzb5fLnR
JXhMNvLWZTgkQ1Vi4m0q7SyzjgXRVu/kU+KpMrJI/NGdEHFZJ/Y1Ph9ny+PpAlVe
n9bAtBQePcqN8ieykBgFT+MBBH8Hx1/sa704h7HIXquxGzqu609gSttoQ1b/t1/g
XLjxYFR+f3tWgIKbTIMD8/c7QcXBu7V6x2trsU8o/418K/9ElD8RRZ8/OuYNBrJi
9pvyko1XcEBMAGlffnYHePXZXpNRBFORte+Hz23uQ1BggakcK/Oo4UUVct1HpGy8
ClwGyxh8rGuhSWZjM96CxwE/f6txaRsoOwJILSrgTIylZ56LyHCUwp4Xjg1y3tDs
O39OhjfWgRLtpMrexPKtMh1wKxDmqgLz93BH1w137azJcT0O7U1QSHCPTafQBRt0
R9f+HR9QjQds7WVk87C9DcBr2uHrYPvdXFafAPSu/G4viTN3OkNzIPIjcLUcl+5/
1PrP4cBDm/A+FWOHF0uxo3AGuOZ2KAMwcHQ6uTpd1s0Fd1df9Zr1rlWnM0xgmY3q
GdqSa8wxBc0om6JPMHBxIS0KKr0TskjDAHAdOGNuHtXOkZRG4+riZrdrO0guU/1p
YWJQBKvU0GpYheTwRP94xQRcgNvBWKEQ7dC+7UqlIiXi1OdcWP7axmdzGR8nKRgp
cGAJcs3l5CyDorEM//uvNeFxFvKXKTPJsyVQfW2diVJMVdpokUWD5iv7LGELzt+d
Gr51Stp2h7Tvmk7Y0GwTXjCY8FlWYkzglDNA3LzIWil72sqzbnr5mXgQHcss7qAh
WUk3CaWskeKzXw1yypuWhD/wudvV17rB2FtGkWSzf2xnTKqLteH/6Q21BLUp4Bdd
VUI1DbDQ6g0gSI5GKiW4hRxGlByV5GVsL44w5zsuZd8GzLtGmgtE2wRJanRz9/xc
ybfmiu2PaTyg8+npl9OvN9NbelZqAf0ZAi2XJceeurR9nYmfiX/hvNYrTuLrE4QP
ppZmVSwtgwfkytjKptEC1Sh/+1jU1qVXPlgHS3QiOH6WvyDiJWo1JyVGw7napHpz
AcThlK3k+M8Ju6b9qwaDRfGcfi/HlbxvDj7hk1JzxYOeUw4CgKTX/uiQVgTFRvH7
sD9riY7CFcXO2Qo20Z1Rftbhv4sCZqFfUPCEotxlo8HT78Uv1ro+3q6K+JsAxaf1
/jB1sUX9c8AimHQ+/Bn6lCDL0H2xEeyDAaFa6Wk45uGY6ycv/FiwttFbUcuzIZyT
uULV/sIo/49DnyJ11wu7/Kv1JRbMqpp/Qhxah+7b9iGgLbMMbMOe040BvTKPIuzk
HsWM6VSmcM9SggS8DkFrF8eG9E3pVFq8/B3GJBAkKsqwkSGvVPXXcs9/mZG8Lu2T
a3I59er7X4+RFP5OCrs2RF1dxcWe7tMkH6lmCz2l1gfTD30grblUi+0akwdWBsip
nR4IwHoe3yVycBkFbDlvqcWq61SsNp9ZJBQuYpQB+0E0NXuO1aYFT1t+kClOeyR2
k5e+skTlnGHxmyCSfltkGJ6cNg5RRHuzEBuKRiSaAsG+ufRlGpq58yc9n9tdLyD5
Dd/mkRSsmTKgqJWmUdKpK4iS/QDpR8GIji2yhAU3joe4tGbL7pdAfTKTtOQbBrG8
/tq/kpvSMIWzz+B6eRCQ63XlzsWuIz1U5ScVSxbVGNHut4OMOPftegp01cjSodMg
r+QIsSWqkM2sWfNGTm9/EWWzMX0AnUflm1VSOKO1baECZhEYVEDvEWw5if3cLfBg
anO5U+5N6VHqTZZ2ElWH1rtCdhJyNkUZLeCSJzg1s79NnggdnM28kXWDexyQUX4q
LyAaTGa96RK4oiMr3WhioBg/ccjFlc1A/tOfGDWGLzHANDjjno4EmhLK0wq6AHg9
IeSasCjI7fRJpkd3FbmXeumlenX6ycvaJYSSiL88qAIj6NW11USI0yAYN5TV3Zy2
bnrcqyU2kkeCfT6Qy0/EWxbaWdVzMYspElSRdNsUvCAUcPBgRGY0GG+XNxqoQDB7
/nB0aCN2erZ1npCP0AsZz6QIKPJ9Ce3wMmC8FvxS5UMODMZzEhc5X10/iSW03V8j
qCfUQaly6zyU8gBGcM40U1/gxTKoj+CjT5DwGG41LctC1YOVNIlqI0Kq9ShVnq50
R1uotBknExHDaCcbyge7XfaUvl6u3Y2Fqg3Rz1424W5EVNoRmxBJA25t75LLVGW1
mi/JqqCD9H95oVAiWwhjTynDVxXYYsqUSBKTZUniM3Rlj5PAlnbn6g3wuTOzkIf0
Bj7TWm+kzrwVnDtgpmVrxnuwfWDjpdM+Lxlxqq7ljCZPgli4XCwSbKctA7+LJvSA
VvQN2z/R+Tep4AfbBEYAjDtpLYmbsSfcVaWWOQiJbJdonrx/YYwyErCU7RxTqdBN
+NBaxqUwzD1xQhNSFsEoDD2S+mYNI5i0jiZcEzkBZiy6SUSRzOjgUgPFMqCfyRpS
3cygIa44eO4NKiMtA2HaFCm00trockvBqVBhiU6P0PynIPE8XaA1mETkFoGOpki4
d8vko0lTTXg80hjP3nzllBcOcTWwE4sTmUbI8fynJumxrq7WEY29LMwFwH+goWht
9e4w8eqkKZtNWR44Fhbru5Q0HlMFBaHTM7x8gMFQZd4f40w8zMlpmN5NjsY6AGGJ
JaFmG59lP9m/TESJ15lpEO7avQ11tftnk5gKQPfwHCh852rdFHr/X5F985H1FkaL
KeoXNYDuRFu217jOBJNg40ovKZyt/pDYko45Ob/sA4mbui1ptF1O/SisdxbfQpq9
1MkF0GbyjsySO90e/nxvmclSiYU2HIJFg+WZCjCpp4gOzzNv/0L/rrRILHu++Zgz
EW/V+uguVb/6DfV7LFObI3uwS1B4O1WkzCUne4XVRQNihtqUi+njQhAIZOcZmg40
bkJlwrC6CsITQ75woDvRsX4ESlWs99fHdV6/OxBD8A5Om2j33/F7EWdvaBU1qCQL
sO8misvwcvu2ACJ1AuuGcb7yJpec7H0/9AhkN9Ai3uUSCbWI+bRpJRu+rXRKP4eb
XYXsnyEBPF4urvcamilKgBmREFsmAQshOttj9TQC4PUcpiGYcSVJZtN96k0dkUy8
RfAA30Y9a/YiS4nowkTjQyYnky+ndaHgjqPPPjv5qo06s/JYp411uMqn5auns/iH
F6VevBn97zK6SZRoH27qasGiSOvN2toAbYfaKsbSKylZDbfWuVOyTtbsbKTI08ww
FP8pIRn2qK4ZLNnegf8KvkIQ8ZNOoODwm5fDPMHJipzBxZV1hAcId22x+tcyq/3d
ZvCvaC+1nyPNafCRA4grFe4bBMPsWkOTIXqssbL4ST6CfBvS1poF1pyG30A8uKZY
1+cSAWeoEN/2OTQGsz3GcnM51ASRjXSLLNhvwZKawdkj4r5SbDSvlCzUMyBWNOOk
nw3IAkdZhBgzV63M8ywgUEhIYwTOaAiIVP2LNaNR54/ybIYjniuOK7G2MCDH+pUb
mUpgb9gsisgZrVFfgt5Zr5N0HASd2GfEDq81t7+BDGgqUVfvKNupAFr9KZWBujH2
OoR8MVW6ctP2RMcD57lV8LCXlf5U66ZGzHb8bGI9WUTiZjrDnmDX/420ftebSxF2
fyz0JNbE9HNjRfupFPtSWEvUmqXjcspMWTtlMAkUkn2ipskQ8R09udDZ7CCiqR5T
WJ387oqhoCD/d38sa6HjwZY4hpY7zpkWhGhRpWpGv4zv/fDFsXL8bSTDqsCGKti9
eE9ab6+fbulckaC/24tKsY26OW2ZTrQzdwQSwh4UeNU/yz8oYIPGt8VnCRYBfjlB
6gzGlFPEw6u3OiFAmvzRHUhdL5GWuQK+mcyVOkuCX/e/2K0RsaY0c+NgjFmzQzPv
om1bdZ3kf90C7eEu5FLx5TOHUYGfZ9jmabnsk2RwRim5e7TwYM1n1Sun1X5goZWb
4biObSZCqIosbHnTIqlkgcAWHoygiexhfK9DkHJNzyiqc+OjYgDdpKvMjCbz+ZAY
yYHBaDxC2PuY2r+6QYkNVC1+EdAXsoesoCpQ/ukVZ1ozt8TSZVO1q85uMWsSf4WW
BkgMNcX2y5HHGVENOEoze5aQJoF0vmCzcVaEQcMHRggj9GtHos1YCAbLTNKUSKa+
rsKBcuxjNtVgoOgu0a26K805NGR+Yhgymxl1afZrdUp+6KI6XE1aujiJvfMMIpEo
wbzu8wAX5qTrWAxaJv4WR/y7AWkHyLLSiYkNtqDcs1mHoaZlpCzbYCqDNgPc/964
gQBX1CSkMbVSnN2DBRRKMVmjKAO+/XNikbT1pzM2TVgvUlRaqZzBw3/V1LxDjyAN
UCPUfoRJNJaKwTGw/pP1z78UOVW7bGYWrVfCOGP78Pwchj8MaKutfxGavbhDq6dj
ppC0coD+sd2GnSgReBQAxW4TflvDy7joLhb1QYbRN4nZsnirDo8f+sI426qjClSA
2QX0YWHHN1Y9B9TYPiBuo8YqRSPf+PLWPr6pARz1z5UmcO2YmWzqw3K300p81vDY
VvgWcZhAcG0TcGXSVM22HHOEd6mTT4DTYcL/yzl3CDg7Xj2wkU88CVlhm6qiT2fT
2o2eibIaiduxrc9/9v0VFkOvWPt06AEH3ZnbNBex5nyHA7sH8o5nnTTj7jbs8F8s
dx0QrxP7+DGR3Aa6WGZkfE7FBc3SfUfHjXzVsGv0s+UBVQ+EDe1ASyLsZ5wF0bW1
oshajpBdjiQAfm+VZHL7aO4Ckj1Xz/1Omq3MYWOaUQo1R+scp/DvWH2+kiuoIxhB
HmJ7okdvnWLbblDgKm2DXw9Z18pxf7t83YVUP9jhrkEKB2QlVJew1sT5IBcQ+ZaQ
uJJQxppJerSvAMq6X7Beot+Ub9ULQ7xjIEKOyfVxLwx8Wt4IjyfIE2vsmv541OR3
z5JlKT2285jUwcob6NOKtqEEo5qWf03FGzzL3wRdemIae3VkhBMl6qDrRdekbP8M
i23bA6vfWc4Y92fDQKf7TOUG8XdCQm0W1MzzoTwEX7DMwKO42yIHNbHDvscNZ9vl
o5LU6SCFPr5g4r3k5RfgL8q/Borq42aJt64ctq0T8vQxfWiYidZXkcPXHVD1BOjt
xP7iarn/QX5lDITrp5GiYjc58xoE+/E/UTutzCpoLuuBHFb5UBrSkY7zqDTO3j2v
N1mSZaReA491GJqkwFWEPwPSZalDBenLsXpCBGzG0enQSKAZsNoMyUTJBoZ8UvW4
QPhsSgufaBrfkLOW/a7LPmW0bkkMK2+GgpFUieKsOOHiW/OB+TScIbZtvBpmfCkw
aa2PQtQc8dZeQtISKXl+IPUm3eQRyiJAWhms7gW5QH0hyr9d7VP5ffctOhF/+6fH
bUmXP9cbS0MBqgqB14jUpQqSDnqccE3ANfrR3ot3/3cFvd4Ndwyr7t/8ndJVrEFE
o2lZJE/6EnoXqRvlCFm99xe3rCPOPP4suseBZGG3P3ud82FnUaH60Q++DTR4DOX8
7H5UAGNg1MBBNcnu0D+8eH1HVosjP/siV6hiQj30wRLtWhaj/VU3Vd+CuVO4bu8i
Z3M8dutlHR28RX16MisWhq2z8t6y32vCacfA/ugFdr+79Xqin6ekQvsBAAI8ORMj
CYyQDzbHFFzxZRZQSma6CC5gyfVWHI2DHi2UlzlFWGhpBqmLmENz+XS4H+8TtNcP
DHgXkuszWcS/2Qds6xLdvW5qUlvH83nXyjpWgg4uR0M6Yu58WRNc/qt8gy0y4Cdt
peVY2R5BHZ1G6hu6pxgqLo5XKwR62YZYpb/8exnsgVjx206L7s409WvcRKzC2+kc
ghRXX8V4W1ggjjBb43pFfjLrfIeqcXo/h6R8DZ3JAnaNHCRrAbq2/GAT1UhlPTtw
tfCLDcsrAhZEKTJttmX0SkHiFVTRVJzG4bpFsloD5fiKL6Ox1sIJ2wmGAyE1OFt2
qA0F4VxT4CSlQqH7ZlVy/fZnr7l9VLLXY6Sh/NVPee97S1XYLr9blXlp5S2i9N+W
/RJH/D9PqNr7f0pmIUVg8Mk2N32jEEbC8EAhplNBF7swTkWRNXS1HlXUMcBuzaBY
UaO90vj0HiayEhlxBaZywmzKx3h/2EBxD+XL4kCkjZj66L9dOkBZ/i8KdpmExHnR
5eY1Wbl9Xe7EYk0YmFvAMCU+OHM1hpE4EzleChbLkyOl16ov6L1gwqTR5J9QcfEz
lH5ZbvqhVVH74p2C+9QY3YtYv31Muu/0l0DyZk+V5wSqMQR+C2fjtbzAGHBEPmvE
509AssSzgdG3waFxgWHDyFZU8pech3G5LkWmhxhaW/Z8FCJnhfJBaBtpXXk5mbvs
HwyJcZ0R/vXgO+b+nfUqJ/q0RKTDxzTaJugooyS7DH1furI9SipEKkuTsSsCgHvQ
A0FEXHNZ3ejxvG4pEPFprXzz+qvZqYCHgzk2wZC6/FoA3O4ZafHH0VKkInYo6Ogg
hpqY1AqQhWm6F41yMsXWHR1kVx4N9MzoJHr/sfItMqq2cJ28pKGLgX/gZbPVTMvH
Sfc/sOPyZfTKk49YfP2w/ZWM8DpunqgCrRKBY9zSSgcKdTlBIc/BrJIm5eYjo33g
ZM6rqEPQpizj7Cps3PfB3XvAtLa5rHwehYjjUfZiJbTvtu12dKd+7rfuzw8sLl+B
Exvxss7sphQJPwjh1K83OXrx3t9J6asPQ/GdLvIeWfUa6LXHtnbbFfYJDDm8DQF9
LEKgIEPST0dMDjD99woz6QUjxt2jXYWDWnDIVmk64wBLSgSOBcE9EO4MSQYg/rJQ
NIlzNmXAyQlJO+7MRjdU78+XAa/v8MbQn9lpFR6bUK4pCvuIj2aXyT9Fr9f5jvYG
rPsciPzg8ARStfGuvL/AtgYcAxK1Ak9gb0U1GFaa231sqpjZaUPQ0w+dTvAMDvs6
cjiArofGYI/WBoko2Yd3obuRNGGyJGxDkt6hOvWYBHSIGPi+etrVmDRc6TYMdSyj
habY511GGg7DKuS7raGNc80Fhy7LflzXiWZVS24Fa1VJDnISgogj9AI0GwSa/cLm
9Y+xee1xwOA9lzzV6STSvm8wPNa0RLsP3OWgj6BNMQ934YVJXYkVAG9cykFpPlR9
IZ3rBOjM7nuVyt6RmF2N0j9tTDV8h2fQ4C+fM+RVgjw5RO3TqrZM+apzQ0F9/nwn
8hj+wk6KtCtUkjJoZWf9FOktT3lsB7CBQ/+aLbbZ6RJoI3RCuy2wcfVM9FuO7gND
gmSnFKQd0v8H8zP4Fzo6Nl6IA8tjaydv9jM5AeL3EAA8l53xQHarxRx2Wo7dxGSG
j3Rv7OfffhfUmxa3IrDY6ixA2HUGZKjBj/mAj4E6MW83SIWPx6A4rNpwMLwCJoYg
WIWI3rNqJ4I69j+KnQnY6h0zOBZQMsVC7Kc1BUBChTHDZqU/6e4gdQQidbGDiz4D
q9G5NrwKCuWjkt4QicdOXkksspvcm0ihYwW0hOTg0tQzm4CMS4YEiWvcskTUOzHW
EFZCpYwDWsSulz9qyFkMmV9qvjKBpvEPIRx6QR+G1CnL3zbakFbGvqOh4WJT2Mf7
Rzf25prDwDKG9GOL4wRvTPavNNHKYmbZX0lc7DtVyB0Eu0fPfdVfrrsxtmVBj8vE
+KNGWV5Z2W1JPgH4eF0u/yQFjJuDh6teKPrN2DtoKlal2BRGQucRinpb4kcWLh8i
Xp5/jKjbUprH39GLG5/i95X2y8OEnYK+a9LVkMO+NXH4VKHRnLDiw06eyt9Y47pr
tydN+kq6sQErSHc/+O4S1tDQIYHUX0ca6qwFoKUHVY4qUow9ftstmNe4QjrGkm0M
QKVwrpUIIy5Zc+OpPTVtR2AvDacobGW1LRSzj4krzEsfQQOuxEFWs8v1luCiqT7+
Le6pUF8flHLyvT9i8LnE7E9dAkXGnMYnhc2HU8NIwO3fAU7ZGZ2Jb1ONHrz4cOoA
MXkjEH7/cI+ME5zNrGIXW3pmcFcAcoukq9ikcBzmQOWubXd2/wS6cevMnfq5rdjD
9TAVjN5Yd/rjLYkR+xjtxnTzxLoPGNbTq3rCvyYVI2meZXQt5gBza0xVLl2bl6VF
6HK5zq3ooVmn8vRdJDGvwCO9Q6J2Lk7Hcu3UWPgRt4TL/D6NssAWdGs7JTbOeSed
rZDm2HgQYLoc8twZKSCqMHg+OmBO+FbX/hq0a+5FkZ9xnj34wjvMo1aA0Hwct083
yqtI8BqeJpF0kmvZPZeroJBtAK8R74gfbe512RJ4+sYkX8QuFLKxUviJHRSRcl7W
tjqOt5zKoEG21vX9BJkC6E1gtLafm/F3JKRCO0Xt+XmZ5T3FyVL3jrriKOZzKRTd
g2df3MiecDbP7aiGXD9u4dVFFeZ5wi9FScQXXcB3EPIZkLf8FY4LtvbYy31JIT1f
MRPNYWbOfdbc0BlowpOQO8h+XLvYqO2Er0K24cb1HdgZJdZtI3aBycBibSVdqH69
YR6c06BWzaq0KsPlL5J3uYgsVatr/6VhW62ZDg8VTm8mWGA5aZXStCI28WllUUkn
U2ZH9gBUcj9TQJRdHsSv0RaAcRmY9zcAQP622VejneAn8Z9vYY1wo3jK371hdMnj
5HRn+oCILWh/GFlLalMbzeFaCtt2zyprGXLetpHfs+d1IT0fI1Di85+BkFpjAnvm
wWf9GQicJoz+CwBlzTsgFTaoyxsPTEiF6h2CSyiclpE1jObr/6bu4dYSzjpOBl1Y
H5FGN5olfCvhZ45sfv6zAIRKnShGTfUSzmpgPTihGyXha+PicSrvMmqq3mNGqwAR
YzZY5v+BiwSBhgu3CVf2UZURc32KockxMMHmyYLLBKo/pWuyQZdvYm7+kH/5snIB
6a+aq5RqU6n9CU8rrk2/ngr9PUFB/AVO4c5c/ah9zoXJXq5za3S0pEQzw30dLpQk
ZsPsNcQFBi0j2Unrk/+8hOSLY8dO/ojCwPIsLv1q8Ie2dO0nwAiFoxVxRLwIrLtA
tI5ZXQsMQ3pPri1MCrzflMs54CGIeID0OC0uPK2X6hKGyut++P2RqAIV2AeKZz7u
LTYuO4myvy1DljgkW3mHJxFlmFZrefmuBOgigZPzEyXTCV+vuz+Dd9ZvWfK1Ht+L
dYvMI0sGoW80+et4yxg0MTa/ymrErNN+v7gpQm+NAJjCKc6Cewx7UOFVjND3buGI
UqyXovmRRrhWPhQFCDq0dFZUhfYxQYvAyyxF63LY+U4+4IIuNnpuHCcVwTRLuqsR
o94N5SLp4uLTH0Y1hX+3Tfb2Kbvcu33D8cSBcLNeUldPHr6ZO+F0yJzqgHNYYv78
Yj9CJZuTrsJK55GJzVdoDiBErtdOxChiFAX9zMFtgl6Y68v4yxUcZgZ+Abks7lEz
WL440EDm1mXcCvuHI9Zx0cAM80fOAW0Rosb+SQU6opteMVIld+OC/Q6uJ4uB2vOs
/0pjX97s4eyzOIqF8iM9NLxkl/8ECRLFf8nB/6hUQkVV+mOEo0qhBtKf3WPC+Zmc
VKGSApJdhEYgQr1yxVAOBNO3GMigos4Qb546D2s4YmnOgMeDrUKZu38lsLF2yZrh
6fSHC9GVT2fmNbH1UXuwX8ib1Quz9fwAiYrR+JxJWnrXans/lb94Jken3JHZIKow
b8oBGHRD5EIKgvmmFJBB/RWkXnONkuchlnLIdPoMWPlc+3wMN8Z+LIYSLeYjVueB
/lcGA57JRKGd9tj1QPJx5RsW0lQQCIja2vdO8vwSBy6yq6Vtju37IVgCBejyHRV+
PNpQIB7TcninUzBP5NQtuiJ1hK7E6SwlAwhNsOjNj0X18fZXjsEU7/cq8+/9EKh4
Fd745v2HlveSPAbAk5PMM9WzMIfZyn1weyP0PNVP3gxaefHSzJdu2MfhB4RbMAXD
Vb24eo4+ZolvGmwdVWOFLJCU/FUfJc/6AeZvQkntQGMB1/fCAss17iTj3arPCclP
PI2zFh8DECGH0qjNi+14NdU/0d1yG5IFG0MUGEeuWop3PmLq1rD5QKxU/ZFfcAp5
V94fSoLp6RL0tAsEAPk0t0heJKE6nLdt5gELGWq4K4SL62Y9U5VihAv2oiuwANVZ
RaYxq/qwg32OcQBt7a01SJiJWf6vBGeDjOAx9HmAuG13nsC5Sx/o/aFn+L4jYHqI
eUWS/EC4g3ukbwIlkcKRKTP8qmv2rEt5RnNBz054kG9Tt8qfq27ddpOeOlcxfuvZ
zB8xj+vQl5eo6bKJhwSGwWTipp0d23W24FRu7qkURybfgSiNYb5Q/jKxegTelbTU
0MC/s3oU3DFwt671+1ZYsGA3x1D28MZio8vtbetuZB8CC/pXCriUuv60Qv0Hc33g
XNCUo2dcC7E8S+eziGOiHjjvllD1LIwqa8GOthTNRqeCr0vN7lQIBywDw3ov8GG8
dkI3L1u+zs/LbHShIcxHIO/TqrIqIYc+Nqu6VyVM17vPYDagPZAshBHhxgbeDYY3
gXgNppw6rvUCyThx5w8d0Rq/HX58hn5wCM8twUglCs4eHI1YVsH3KkKze9IPwUu6
r5IogjvD936p2kpG4J+hSEnN8mhp0k+Nfe5dfmZnp03RfevtSqrfF8ipGPE2aRDe
yjyicl2xcy5uqEhDGMVGsMhXbb5uHgaREJUPgFdwM0Te7x7NDRymDV+gYn098wg0
4ib9Zo9CzNIcAsmJALDrMdTeyarlu0HGHHl78PoBPHHIV5HZWU/1RURJyihVeot4
J9SNLM9D8vDdQ5YTkTeKJ8p9TkarFkBfRd0NmmpHYNJV0uovkOI5ZBoLnfpsbS24
OT5KOgdOwcn4p/iSMcCUGvX7XcZG8AX4es55tqRDS25eFDmGbTh6HhxXc4FS4sou
ejpdYsGAsbJ1SUrK2Y80CDxkGJKtC0rMo9WI7t0U9/pm0AWKKUaoCNZgzLKbSGfn
FXmnod+A3F1QieDvX5fqV7mDfh67PGOT3KjWuahJrl4VXoDNecq7d0gkCeTZC+Cp
vWPrE8LVC+cBTjEr9H1fXrOVgzyy+LqpSgSzgXQ58NG8QZZNc/pHOLg9IS2q/wV/
ZAb6s5H7hOOIlRnqTbPHs9q7Z2kYlmWgJVNV3SM3+ZFA769PJxdyxmeCmXgqdVBj
5WTHFmvlqGbJPW5768spExdzzYC9eIdEztbrGwPTcbmrtw4FIs71Os0nwkTvXxFU
njdAMVyl1IoSst50b7Qo5AsCp4y/u1o7setHiOQI13krNWzxpXElqubvmbC8fK09
aNPeN8aQw8YHCROo0N2cRRKBW+UsF+OcucR3kPGpwM/Su3aBNsRhVOXF4HcjCyp5
W3VDYzoyLjd+U1VzO17pmQHR+QIe30sM1os9/iT3D9r5Os6J7t6pDVzeOzytcTmJ
SSJ7dupFMeygN2pXqCXLnuPNBFETdqUDlJik4oO627c1dW5WMs8aQTnqE8QkCHvI
ty2DzY9Gso88xXTZnfZmPKTbeTUZHL6e1nCM4r0xByzveJprpbwcgMrFro4IyiKs
kS1NoVNDhGJtPoYoVdjwXzkOcD077cZdfXjDdZnCATL8qEwfd4//V0GMH5Gsmeed
WBbX5/nW1jHsw4X5rOpTveB/DxmWM8DigVJgIgNg1iqV/T+YWoldq2vkV1cDKcq3
80xTx0twLmylgqmSnVn6YMVtVvAU8yB4rzCXA7Xw7puL04gDV2iMeoAdSUxxUKFJ
xhtZ18LpN3/Wp+AbW3ELSJ5VzUK22MfUexHOVTXQi+mzBVQbgZHEOXwhFYBjitlp
1ToIezQiV5uxwRYA9bWkZYDJSWNedJOyBw/pmtOh1IPB/Ev3t4CunX9ME71HOAtF
wnO/y+5Qi1+Xr4s+YDBbonwQL2asjytX0QEA/tkODf8Rxgl5+Q8YNoozjxKAhl4J
M2YYFyHlsZViGZYfbsbowTS96RasTf7W6UlNv4O5Uw0QCzeYvI5VgFijHEmRmAVn
GXp4B0qBtEfzyznrvjnXOjiV2s1rQEomhgzQrFmvvC/KJzGjn51VND2IPZuhnsz8
9QzHRxxiG0gL17ByjGeGHNxIpUb7jmp99KuBxyy4bqupxC3iJnropZ7vaa2OICj8
gqobYVtmwCkOWiIZFv8rNQUdV5AsXhWdLf1gK2dFUlvE25QAjc1FddKHwxSIzQIE
AnUFgwbPjY/F2OPWgY4izUsiOY2/NtFle/pdAtEY1TfNmtVgusjvx67uwLpo8n+Z
UslNRcDvHUX9qbI6YyMaw9BhBuUrIeGvrBlDZOSOTIJunp1DNBgMd4RdXo9PUGaS
W40hNPVvBU/5F5ABa2vSpmSE3CVbh9RPltPVGtBbNov3Xn2HjjFtwJl8ql3OJlEi
7YshfEhUDbPmZ8VhdLmBUVaFHP+6KbxuCnbyw5Da/YXV+Syfe/hOoYIXGTgl5c7S
jJQFGms0R3afu9skx6/FQQ/Dlu1iaQefXJLvIm9OlQCWXtZccX1/feYIAwkPJ3on
cuYWePp7W48qb2O5vhFofOe367j3okeF//F3knqBBYiRqTzlD0zPxJyUP0WjS+Ab
+UFfKNIHDkbwYarQ/7h4JQKyk8LFI+1zxfmyvE/zZgYOSDSE503cZBwMuHOSNBqN
npM7OrzckByYXqAnqei+CPNfjsdPW8eCzyrV+W8GJGfnofkuTm2lt52PJ0kkUarQ
NsV3fjY2JMiA6TfILBF9wejunHPrY+FGrInLgpnr/004zEf7Gw3dkODAzfGzoxQ7
Xy9LHdEpgdYu4zvI0CXTNyYPa253VSoj6b6Tz9UZqvxZe3RJMq8H92lGtiI9hjcN
zTU1UUEMG7OeNP3Z6Ve/yxM3+RZdri7dkN2+m0m8ns9+PTxaJnIEJBVq3P1FBu8I
o5v8nrFhR5IpCZXbSBZAArklAddShIkFUdXUrpRrwZdbp5qBqGYIVNCU7dGFflT6
ZUSTEg8hL+j675ialRLG8CKIDLKoAJ8DF0711CTkUn3ZqY1P1uAcG9SgSaf4vtz5
wCaidkeLVa2dd96RX91oZcapPlly5hCZMU9sSWRu2bKaDNxwr8OEqt7nQAtl9lRR
bTK7xuJy24UcW2N4lBZ7AcZcJamlCxS5o/Zmk+Tq5P3o4eCpP4D+jHVVtP2g7ITR
VaHAIx8v1+cDTeTEgq0EK8m28iQydtR9MByPTlEpo2mF49fQS+3wxYLYplH4QQnM
Se+b5wtrIWK2isaEezli5coItnxi0gdahoXrNFvFDvPLTVuRmm6m3uRot+tljWRV
u7jI1uZMu+kATa8XUN4O8Ij6Z/tNeuSSJVL5kIpqJ/flq0gqjIKLr8+cVknatZHV
LI+3aMtqaIuOdD9TInItdWr1tF91CGaaYrfJGy3mi+ZYAa/hm9oF96uUFMu2eZsD
xsrDNVoejVnFnjtAzicLTjyw20513yaVdVr3F9hMySJ6ogOSAk3hY14JM4jaFMe1
i1ADXLP0scuzI9jwLmqfuAIJZuuSWb4SClBGUiDmR/Wc9W8Vsyk3K90+ygW8Xf6+
Im7bB+SUV4uhhcbQDJOimwaUVeeQw27m+MaxcgrnKD1nTqsNi6el/UCrPk7zHpYn
r6MPZusE+wlu9vxROhd4T77bZzi7dRirQx5c+agteyRALk5Yy98Fn/m6lbFWVcoE
d6BsjVdxlvIwyczDRpg78IcYGsvBPaeZyiTCo+ZuVUz57LmhyAKct9iYJ06j9Uio
j1JXB6o3I1caTOCtqRUJJewgL44jkTsh0esk9E8/yjQOboEx+QJF4Q3VwEnEKYIm
KICxVXL0fvQKcVZPulHC6GrJ0AZ2DU+zq41+LyCMCAAtMQcyux9TvT4IKqsabbZ6
iLF2+X2OiFvHfLu3kOTHraaI/usJoOR9e2kdwgs0stRIMrdT0TqrBf+NLOAC0esn
2ZNpwTOwT5kSbuK196Nm9UoOlGY6U6jlxlS+WT1dvei3qG8bnCEINIOCDlqxh0Wp
ezUvNeSfpqQ1S6hhuQ/kLBhTbN/Qen13OuHbzE+YDTptKhcZbUI8j9+wWPxc8+jF
hHQV5AA9S673WQSrYBfjS2Khdry5kLe3CCqPbBlNTwtJStmAFTi6jDTt5IjUKIjt
Fqf5ywDwwrKPFglVebXdorgjxyiJtdJL842dLWQmcWbMIVonM2k65tF3C0NY9K/w
3tGAGbjcsn0wrfo1wUyihESA0qHf5ow7CoztXBMwHZFfA/hEktGDw9cJKbyeZQkN
I6DQTh95RUfcgM6IxHfo7Y/fwmTlL0QCICsRE1nPssiynUqBXlsIQaiDO8+bHO1Q
SIl/RZ3APH3HfD/TY0s9/DbyMd4HGCvOenfZ1MjB+ioC8a2/zQPG4vkndUFYXqAx
ICsu5e1Y0YVA20RLfniz7+tk6Ct2UrZwCRb1fjju1FUX8GOCxZ6/kc/Z/NMZeG83
/RSM/zWCZWrtg5QxpgJp0+Oc2xjj/bhNRi+5J227m+OtTBxpl6c5S0LESczlymjP
GRdspgzQydZGdKdbLhZajE73hFaXFPrb9BmuCbyMYCTEoGYqcN2Hu5lnB0CJvV9j
UhHpsovgr4W4ijDcNHnYo8U32WknBttKI5fkKjMmMOaqkTcr23DPLLkV19+q2ZcR
McY5gG+mdmYUR5i4IBpcAc+2HDc0PIlK0UPnnCM8f8mk1dOsajyDSYoxm4VIYJdm
Mevi9RctF/oO0pk3oFVOI5FIsF3/mxgICu4tqn5ZZbOR+IwIW2XcaFsIn/Q9FBv3
RiQ8Zbxw7FSUvHlhKTKZlGyBE583B5thtrhP1qVIGyqbSdbWDmrTbMcajx/sXKz1
ef7CPqdH3QiKo9/ohjbWaIfoMCmRM0CxMz/bBwSGPKn97+bjuZNDndxzdEF8I5s1
+SzDSXDBYHbF17TAsdiRAV+MmZOKzj1otaAEX4g4cDVnxtt5kOBo9MU1k8NOG1Oy
cSdryDfveuzjXnpch7oQ/tsjW7OgPkA8XnTD2qAFg7RmAHQshVm3Bti8gFdgtl7T
ZU9yhToMBNIn7QTOUdbKyDHrRP1gzp1CdQGKWeW2NA7Xzx1sdEXOez5Uwjuwml5d
6XpCS73213ZoJy9alJhWmiqm7XmnbJ7Jj0nRzTINKD1R15EhmF6HK8oypTiX1ciM
miPyxvkEMht5r3u3vRnv9zlEd/G/xl1qxtK/jcmOOldMDMu0q4Bbm2tZC4HnExFX
r+KTFKxqm+sFW8zFDq0RDEQBgw9pmRkPUN379Gaj2WCPmWGuSa/g8UoeriZ8/0T/
QRWZ020FdsbELNei2cJZtS3okOht5hIGTVqMkUXffMDITjJkxhwwCOZaPPU0IOmB
IsEEyRq1tL3WqtuDFNdpKT7EOdq8P95WFwHXS9mXfnGs0zxAzEOdR9TITwkeIihc
OHkhkVLattdwNZg5oPcVCmKBfA5hSz8ay+VcFutU26/gGPk7DQvRmJ4yxUFwdDA6
ydhztOWwTQzizUlCkVRDqNG/rsmo1JIX1lw8rozJvIuIihcZclLw1v1+XeF2G6df
lskdwI/ZO7OHW1XdJu1OSz4DBbyNP+3Dox3W5j68vnr3BWuEhIVKAXA+tYLC3Vmz
BR9YaX6nTutHOIzaRC4QCiii1QzUXk16Wy9x0KD668vQ2cDXoozZqJzD7HOHykym
rA2Y2HcVrC/A/MhIvUEZzhAxrp/+5qvgYF9a23KhUNUSok8EFBsiLtGznodg13xd
KHbun4aBulB6Qw9BJTJwM4IoC5w2i2tAM1fxAqHwlrzJrxSPPNDT3fteCwmumxTr
E1N/+AZagurJk+wLoV9x60WTVQYw1LxSIGwzVkxmoosVeIrXp7Y89TGs0du1hL/4
2palEjGJgagR7tdnpCooFOOK9ZoCCQvhVHueYC6zgoNofNek2gTc9HvExPdUbGgR
RNPoZpyU54qpLy6INPwUXLT2kzc8Qdh6NfNpJBONuWuEgO7mAVBPynHnmh01FOsB
WHqZ8gulOvIGCkpB3l6xw3e4Ry3iudFN0EW34PcQNsN/NY2CWwqRjClOqcYxwojc
8jEcV5gEdBrQfmZH8AntDU3AM1/LtgMxye2t4LS53sezpdG/P62bFBZbgUGoox3v
kN2a2aWdQT4HqJWVdh9nAdTE+i5TGXa9LeBW5GoPLRVXvXHCV5XY8luJcxpUghyh
KzXKQ/NbNue8w7m6ufcCMiCq9f88GEHaXyHnYWbdfqrC515ypklj279p+G3SshIx
sOPpQJkFIQhOLKWi8d9OYLOzMfep0DbSOoTXTRpUOXlOSig4PmeFcorLBfdxNuA7
ZxH83QjIf0gegu3IAow/hKi9sxRmMM8wf/uzrvLYzB/qO991utR+zIgwQhLNflMb
TPlesZc6zjwgMYn23kxHekLo8ncjGS1+NMUtUzRzO/KKng/gGNGvvRuU7xKEj19W
xnXcTGJv0ikQEmAM4/Y5LQtkEjwW+X9jbYKhsEcgrx4xvI13BUlODNvS0Nqi6Jkg
oPlEn5Mylwh0z0wGzovaThqfD3UvUDVjf7FHVM/iYUwVgL12BCJCroZ+zNclCXrZ
s/LeC3LborxQDxVHkkZ8era27lOMJ3MRXr1M3yvU69toZxmVo75zyPa0Fr4eg8JW
A1D2yI3VaO8UYh9IITZQEr0MyCHxOkx/LEChSHNtNIaG6cnWhtZSeiaBlM7qXs+W
gbZvfLu0rYZKmfFrmkWTvceOIIoyR7UI1nSGUwcjvVtynHllpycXd58XVrqe+lRT
89IL4Wjiu+Wh/uZ4jwbrdShcqczC1sz45fWVDHTLP3STwj2bca9dRiR35MjPmJYg
IsuOsWfNFHixcNAkfdzd8+6hSiVqfdUwLac8cu3sNTfNqJynLvJTYxi6V5ZmyhEC
oaIKckoY0vh5YWgrsC6fqXT0svUCemVt8tv5rjxlOai4mZFhYHMRNdK9JdsswMce
r4PTpIv51AnJsbZLnhamE8LEI0QL5uTUCjQ1CG3eXfvkVU1+h8MpDoe9CF11Pe/S
/dHlfj1ZrUSgS2JTwtvL3ciTcBxVr4rjyoJxlq0rN+FK+zkDX1WP1No28vEu99dF
7Z+20ZFoiWgScC1wnDU3T0KCtCvVwi1oshiUNCfAOTc8xABLkG7b/wjqo3NF1V1I
ug68SXubPZiZSnc4laD4cCGOb3bTu87qLLpSo3jgSwswq3CCVOvanMUWCXc0Qify
6vqOs6W7tnYsf6E4VXmX4TCjNRz6YU516M3lbhAJMQNwnWXPxEnMGNGgag6kcSH9
D5bKeLAXldSUbTFXIHzuB7AFQInSWp8bOMhyP7yXQs1n5e7bDiqjQvagHTRBcPee
/cy9v99a5vax9jAcPN1yQLG03vPVpIjy7Nk7bYR4IF5XS87FfL2+VWVePNX2G+fn
CCcyVlAXnWCxpRW3IjU1Zz9+cgoUcOWx5Re4d/eHFi8hkDntmlkrzTdviJP079HR
hQYFIO0MmP837XzQ/3ngL+bXRAzYoIMIX64/0UMUjOlDsJ3aeCZqcN09qvRJ+dWd
lxaHiAP8eC+FutrUp071bcai9z+4AiYW24ESvfrb47TyfjBQ+YTyyZqtnCcZGnfr
XYzXYzyo2t3r9UdPGTZ4nFoydUvsd8BrP84pNmNr/ZhYi2LhEn0k8RAKgBH5swpy
amsH6C2QW1lokA/jI+RF7FB3ZaMOyBe4grfTywa/AgwL5EnsksoSn9ma0jPHv9E6
wSJd2N1ivNPd9r36CpU8xGfmeZidAl6oJPK0/NqRRdC0OKI7taXXkylB1FKYLGHa
HDW6MQ3NXx1XkzF5ZOGD9rDriu1S1FzW8WbqBVLWIF7NcrR5LnKz2UsW9INVbKkZ
wWBh18ZdSiMQZL10aFD2ZT5py1OVa2IK3eCJ01le2F1a56juDNsI81+YENY5dD2s
EeTnt0f4YiMlD99JJaNqF2LLbTeIrcu56NLLU2WAyn03vY1Lgb5zuYMtOG4t0Y2p
5zOW0rybXi8HcFzI0I0CRSfM7CwA50FiU6Efic65kahGUEAbKGQ2IxVrHr0uqbMu
WMbbgnP6nvjAEQ2JWW7zsf/QEVVRlCa490WiFe9M+DTYzh1J1CWcMDWFPuIkyDnA
6bbtt9NY/npINWY8brgifDJzQfg9a0hb5w+bOl1eodaTfTpZeBVekKmnH0Kp0egW
S+WYU8QlaCPaNt4AWN3f+2eV69BHwFz19RlhuRAD6hYm90IitR1TOqEbWX39FazF
oV3LDD6Eo4WUF4mgjGG2awUq3RUuCIHTRhYowLsFc6hCGPhm+y2hWAVwCTmcnvem
GpKK6UZtUOsPuTe5wqM5p06BZzUT6jd/AB+lQVwEA6FEF/FRdPWsIFbTfjcudVWm
ZUtDKDIJexm9tszKRWOtvNLnX/uc0TI6NBynSa7e1psmESLwSaZntsx4MkZNg5Lo
FraEnDypqKkrJj+43yXeLAmrVQpn37V9l6cyxTWtr+ItCPAZHdyoSARyW+k7O+3m
DSBmn7YLDN7e9bmja68JX8tDdXrJCV6U3M9ygFO2YjbhFxJmhkFUOGE4b54P8fk3
9VWOrCNchcEUey6lxct4selkhpKkBSkuHNw54ET7p0MD8jGfo4VH2+uwHxtI6u4r
uFyxrB3iKOlhbwHiUjG4Fr5VAZ89P7fAfCODaczKJUvZuRQG/luVzMTCs14jBAM0
FVIhCmCJe7WF+vz1nc9AxixybKXoiGFmy0qIuv62b1caxky/WjyA+fmd8D2qq/Hu
QaiMFsLsaNk6LHuh1cbn/kMOyXoHRKuFo0kM3bzZlueAYHN0GR/sPCRurzHb2zFs
U5QgH3jLD0zd6FmJW59HPpz59KZ0hiSIrxfE3zTfQMp49tA9eyQMCjl8KmBFeN3g
tj6BmyL0th0dZwol84cR+4KrwBVMhgCg143fNjPpVTxMnqCpEiZOXL3mv1w9gWu2
9mjpBPaEU0PvFEn9IthBxkpQeVypz3qmnh38Ji4iwpitkmuaLeOw4hAb0RTGCd9Q
O3/IVt6laCpv7QgoAMeKBvQ9OGPF4VuboQSb9Gw5DqlA0qSM0nN/GuAsLuUCQ5xJ
GzoHa7zSCZ8QRLzGHNKxkssEnin423YJNJhHheWoXtGUPTHd8NmDbh4c8Mvmae+a
2uZALzGqNkC4m+nnnIG4wPQ2h7yyjj3VHkzBMN8ld3LWlRScZxmul2ndvHkisRxT
7uAcVd/iS0TGOq6Irg0EUOorp2QyWc60xqSLvfx1K3ONgJbl6qQaJQnKqq5u9RYQ
Dk1AGQ+hKFBoBcDtx4BoZteIsCPh3QRei3dGcAhgX9e/M3GN8IVr1NiriKNw7sOI
OH1zbLZm91ibAra3FcO/4o0AAucTHPXs29+SAorI/IBR15TNccqDeHkG457QoUVl
tex0ydESIUUPWV2k9UEz8HbM1afbcLY0R7JTyom2W/enxTNZ5d0zNfWb65J4F2ny
4Hk5K+iQWrIabs40U+ntiaHVP4pQyPBf3vwW7iIdCXtY1d4P7w8u/l7IvaLdIYo9
b4uXUv24L61PzoNRNC8iKk/+xdv8hpyaweP6uvPq2nMHrwKtUoReMnx3JYH6otmn
0f73+CGNolxuEgNvMhrlQqL26kDmU7DBRgqyubj7QOvLCIeFggG0Pfm8J3kBYcmm
Ukd6AaM0MavSmU78iIeaDsKmOcEZcITEx8Z3tgOMLtYzOj3GmOsSdAvAjMnx2+Gd
4bXVwuiYiOLmnp3PBpJPTkVtFpMhCk2ils2SFhD4DUIMN0c/M1c4rouLIcDYNd+P
Myz0ILJ6Z411Hr9INBOi6OepzqigUs677l1oBQHB/41TiyHZWTy0hVIL7dJ/1TXs
bE4A+cLlKSjk/ZZSDDFBMB8xPM8NmfRwtx9JGGgAwjXgkkIy7VtczAjuxwcS38YL
e4zNyQpeKWpZNO6CUpFk+jnGlyW0QdlN/97uXkvyCjY/we62uISfiz0oY8ARku7j
hXBJk9A733/eACwcS+z6oiHGFYv8TfPaP/JbVkFG/Z7GATiLb+7lx5Wnh9rAUeNW
/3aZ2eoVb6MTLruaehbavcHaxpfsdA0BpkupMAN1jDVqmN/W+UUn5v3aGNSmrE1L
KjHY39WRWWzskfoxT3WkmgWbz+oN+2+4Mod0JsGldTMJpemmNMI2r6ozv0sM5BVl
RyVvn92ggzoqfuMIZtiwl+461X6F1KeBq5lDnTa3ahMlbHi4p0fc2wfGxrPBApiH
dmlCEGJfQUrqmXRvt+rc0S5O7fWFbmGhJQ2u57bXyjalPMpI4PJVuFYTmT7TXR66
9Qr0VO0F7bx6J5ddzxmdjdC81IUucSKFsFCLnsXRvMW7jHkLQdn7PLDZdgrZGAOx
U1dkIEP88ZAE234NR+dskwfxz3uPZMFsZLDbnphUOulIjRnj89YuZFRPhPuVqQsH
OL85+xJ0QxgoUQEI6uXJxmcKZ8CYFkiVjCQYNMgmmKjEhm+FPFo0Y4pFu7lYusxF
40ACj+bOwAkBB/+x2qqvopYqilml+w2X5hNcH7Ck185DLiPIGJUVv9BVIjoSZ6T7
lhOJ8ce4Gr3F0gKo1LmEtMHpiem/H2opRSEqxDp0sJY70fZ5uqFQDm0MbQrwsZG6
z/dUdJ/X83RDaiI3dr95pD5qH9AjxroTmDsCXvvCZZik9n9ENbPHO/PgA2TtF/55
iiCOPMj262KMKCliMu84WccsTtJnVci2HQgDY/Ac+jlKxvTBP/31gLaDc/gmVOxe
jNJOQaqn11f3L8JlGhAldS7Ja8XeYepSRF+YaE+DndPQfzb16dlfU4fGeqosfvXL
n9HyZL+C8dSMHtt6q4SSwFIM8DLzCWAcLVIkPPBSZJoLxdRJ9r/5ut1VtpNp4/UT
P2XrkjJ0iCPwOzTAMe+J7SVZVMLWr8fTf8uTNHQJN6hGTgplo2bU2hfKvRAre8Yd
NM+iwIBcXSZ2SHm2lltmELjdf+UY9xGOHGHVkWaQ4k5KZxOPs5dQdkGOEfMoRLRB
JN63FYvOptYuq4BcepQz7voQerCNCFC94pgbJJoyflN96E4QkXRyB1DHD2T7NIgs
l6eWRVAgM8u5fn+ZnDE2TY+KPCq/lgocC+hAopcjA0lXiX94tp2oiqC/0gbJmHIU
c+tHe1XdwTyIczIdz0Ca2nnVjLXkDk3StwMq0ehfN7LLm1Uf+lL5RMLiuSghrquV
JShjxWmaxnGJZy0UodjS5JjZ3dFbaFmk5yrdVxzZFEHbfYI56z1m1QekiT1NkB52
nkJu8wztTJxqq4IFR84L/2HNK/Ge9yhXyRd0WGvCSbtx0dPNuG0cMpSUBYazW272
81X2ZlInPc0rvs+I08ujVfovJZ6/kcHsL4mmOMBAIw+ctOw2ML1OrSKiScFaLZS0
lAY1LDYMO4qnBbDmo0iUIY3H7rIbBMMJ29YbVH+WHnK5YBVxKbYZekrkvfX4NY5p
r3loei8ntiDZn7Pl5hlDc91eEsZMnEy1V8aVQ6ZPEULZTeaGx3E54Gn9jSugKQVk
uDu25zQ6hF459xzxSJTLXcqX1vAnUlwoUs9u/khlRrTuZDqIhRcnXDUmnLXfc8CO
WLGGNyysq6eXd3LZnGbIxe8McONBAUqkwF4wnVEPsU2LjAXduT264tnCt81wAV2h
jXdMclbqy3glh6t7tz4Xs1n1b4yPUp0Cs1xGQExkrM5I0La31whFQQLg4uDYxsJT
7GT8zeRdYEOn7cY7lNnEe9yt87i/HjAqsKDBGU5oEWRFTVb4XiWsYh47srxG7uXB
ECWJ0q6KCDozsVVrVVGQaXbhSTU0nZqcH04MrHHKZy1lIUEY/nAQ245JWVBRxFZF
z8olV6NZOpJD46PhXaDG1y09aZn7DUcsXIzQJnd1rn4tVrw4DdQBMIavCUR9bNMl
ng/x0wu7dj3arBDlKFENJZ+veKwBYTRzJE0WgshNEHw7Is0qBMYASVx0ixmu4ICw
gYDduvO0AVH51ANyOw0Jm7eqaq7QH13BR0LR1bEzuA5qBfrv3K4tuxHjDwDsB1XG
oyyMlzDEUybwDY56vFQJoou+OrjfXGtjPHJdFolcgUVLJXHWZ6WLSVOJW2sDCXbP
YpyR6YsbBTH8rxOkudrOV0jQB8gZb4TyZGvVJfsLLIXeXKGLsNg1r6qpKcjb5t05
k4yeY4nOwlTNYFYm2rP5hMp92ICt8qCRmhUnEElQS8Wo6RR3ved1nU4TsN0qq1WS
URIHgCfJbPQulEOFI6AVlJqAV/qnCxKDbnuCPF1roecvd1Q5jVqrR9XYM0nQNdBS
wb8mvia/1BNQCliGGOp141KPO08Qaf4Pdk6TNJWBkc8jyRZki1hcuhB0gBOtG5/X
qupTmA2Npj4Yg5GqMAxlVgCHTpqHLSmNhtPo5jILcufmQWcamFfGoXJ5QwfnhNnN
FWhSvKpxiNI/VWLKQvhiC1fdso1bIttGHMibiUkw09cCqcTihoDu19hltbkrtd1Y
x5V6RZKEiHNy/z/ttLwkt1ZiUTJ+Om0qPl2w1eMDooZusRZn/n0a8jPspH0lDmdz
KSUQLmA4kWsbRcUTdwp2MSiBQaFFlCUJqUW78Y8sOuCBOxCpk8TYXfcg6LLy0BJ3
lY7sfm07aigi+j/BMu8AXxz8YzxlHM2EfnNsmZ9wQKFSrGhpEXaxbYCOyciWMuQV
wMjCgZ3qdX1Kn/6f7NxUXeEHmMtc6e2gTmCkCbbhjY5SNyadNhyb3PkI2ifmsZRx
543GhWmMskidb1kF6qVseXEVoy075y2pqxR7zbQ/6AvfXhrr2bTd/e3U5p/vv1dp
WhsMkzM76v8aW3SdiunwUpfKTJMzZcOoz/Mtqyut+571+8s0Gh+3SyJPgbiEBPt4
aaFpJ3VKfxLg4wKTO04BsvitMKJ8Qe6ncw3aZjeyAqT7oXV//gJla9oFXbY4D633
5y8K8Yhlre/hEwTrLBO8Ei69MBlsFayT2vetek03uXBMvTrZmeXV03eiFxrMzQtg
b2zuvsDsq1xvGUroDvHJNRNM8wvN0soprOiQDObT4LzANbZGofX6fiDWFgixh7G/
D0EmYieOcb5Ahl9mEHEh6LkUbko1gt3YD1BnCeJQ8oSJD2tTuJ5zgxeocPmxpT2J
T8jbJKm7hoUGjlHQ80FpkKXkVIkBgysSfZsRUjaUX1A4oOj4DCaB5zkeyNK8f4ZI
4g8+z5D1NagBGMduMcnEdbOnOI6kgt86vqkfh6gpssJIF04nzLl0FnUMlXtxQVoc
hRAHtlnZ9hmFw8XtIGU1uhHl45bufo3TiL/bIarefG6sP7V2wFMBTklJ9b+Ji9NF
mLX9xsPJtLH2ugjRSU8Qjy+UjK0nft3v7QOJHBDN4cDVll3Ez1vKRM3N7Z7+pVZR
55neR6mp0k+3DvexZKofaM9urJgBMtHo0DWjsISv/D2IOs+KeCq6sCu7EvO9Xq+H
NNR3vbzG6d2cfD8kXfgJsvo5B2pb3+HhSDBJcVK96JB0DiFt7TkTm5e9p93LIoui
2hN7qpz448Ny0rcogHPyQ1ZCji6gsk9CLN/KD/9Zc6mXE8xBdfQtRMbZZBBLOWLU
vBTv6v1KPGkodW4YiUJYEBo2pFvc+DI0tpiWsUh5H4r5xxgDskTK9zocK51c8iFE
1hkW3bvIPgkNXFcgQRfiPkhpmxrCYX6pXEmZDmmzeZ4HeHNazr+wNPBHRn+X1xY0
Gi4PIH1qX8j1UKrOfWj3E/drik1OeG8jJHB2LTYzac3pWKFG+tvbB80OB8IZe14t
vrVA/Q+Vp50Pf3o6CHctprUwUm/xYCfzWl+gJk1vAu8J4vLfPyHy75Cten11aSyS
qqhtGBFjIA8MWuap5njZTYhL69Au3LQUxUfiTf9LZFMZGHOXOYFLoIM3xLtlyy9y
y/dqmgI7r7KiRdviiENdc4VFWrzcbOZH9BS84eKFVSgr6UL6qS2Y18bq5WCCBwEo
81/EFiLcsoHpmnV2ppIlU6ntGrbhWvRS6yq41Ld4POKwdpop/FXomD4j6wxrwFhY
rkmqX7HwnC40MKrWROddgkocIJ8tLNS+jXukzhsJEF3eFMDIR8T2JwPBKXSMxhU1
Oyb5LUUfaPN2pG79w0KHNfm39UglVBtCj/QtbhuiJRv4VM2m6AL6hYJCaO8OxmxO
ljteuVPorivmyPZl9BclOP4HveKt+q5CPDW77x4dDSxpV83aodqEvbjjblDyF2o5
toIm52quHi8/AWN+WTNMq0soRULRSzHWSl+pLFteXaIzvmCM7gJpJs6ODrOin/Cb
kE1qgnzazWTSqQUmeUSRysJHmhfBACKxzoA5MHluXxzmoBcVZhmlO1Db/rK2BP/Y
X1m4F90Q+MGHIF5a3187ejfPu0RNpbAVK+C6R3L5p2itZ+87PwJetRJvenjZqHKN
W5jPoKsQINQDjapw9gpmU41izjz1IwdpxG6lOzem/gucRftzYOo5mgqrqBllXg8M
n7plKqBhcc90/3RDOf5MyfeaVp+WlMogsVKiOf/QVqnCJNY8Jj94d3pbsLi8QvUk
99iGzhCbfMVObB9aipAGRXTaYb3cQe7nNah25r2W1MMbxHENJHg+7iVz8z5StKIP
4cXpHAvRUaOHfNjfqcDibeD35/GBD/0ptAd9jTLVzTpO1nZGYiHxeRax8O+ye5kf
KMl+d3zcQRo6vS0qlnFu26cokXzmIlq9g2B+tOfYnOyWtOA60wMMte07R02lqboD
85+gqReZhUK3XoVbYNNGpCx7R1AZVIiBoM6KxgJYwoIHhfHusvsLU2tjatmcVRgd
+Q9LfCrXFIOpsbpoEmniTEaop9tFyt1c/g8xL9apKhSeBr9ey+qwg9bxcfPkFKqO
9Im6N66Z63yYwPJGONuaU9Kbdx5p9JyIByoEem6BJoowOzU+MPb125HVvlW5x8Ps
ZN8OkpvOPcFpt4rS6rSHyqdzI2BRC5z306ft1Yzy7MieBmNshUqZImz0ZRJJX3CS
vEsmC6gw0hF/ugldiCDObzvF3mCCrRjky8zcVsbwEbTczZcuAs05ED12/Tz0oslT
GhexQVu7yVcw3VwnQxUqwZz+ARSda6st3ykRhhriaPsn5fNNLIC6Ra29TRPvFGOU
5yd15FuwKgp+7Fub79/dkkh75sCjTmTv/TpaddNvvLoGMbOtmmpiEE0+fNMoGTWa
FgcTKVqgrHziDMf4GVyK9IQ2F5drlC3cFrMDnwyetlsSTPOqNzqatbiadVeQPGt6
yiKo+V3Jdca51ipZjveMsbWVGi49JPFkR7fWC1iGSfingKjN8JFkmRY1RrWxuEM1
PKuMlhCtpXZU1C0o/6vyw4Q7GtP7+FIvp9uUWGUfEa2CWM8P4+5RI41tekVNw4l+
kA/o5EYs8f6klpDTPkEjupvHAbp9ETYnqXA3ttC0hcqjt7Za87Er1zgvTW/N5T7t
Lw5/TdmyvFXq3zkMuD9qx7Jg0XQlrTGQ8wN7JiP9xpCbz+Xx9ekJQdkjXRuJPQCh
QU/TzWmp0/9kcXku/ApTjlF5NghSfEvSo+s3PiLTC9AJpftr011V0UWrtXUthVaT
jtMDRJUeMndN6eul/MQlsJ+5klIVR8I4VU6jECpa1HfO27CkuCu0N0LpHP40xLIe
KUQAOGAhwT0R5erJX1kCJXtGuQyMxb3r07Bwy/GEx43tVbD27rGEpuPhMksZPHPL
/BRrDx+W1O8WFMTRGVIWhLcnXnfsh5Fuzlf58dIu1vyESErOvRJVbug1tCc17GDq
4AHxHdvtWmyiXVEfpO1089pbrimrqqxVKr3miNzQEODO5oYOoAJalBJ6ojo9u/Fl
pkclFPGVztVud3JZsfcemJDRio9T2N8vpydAskyVLEdUblpH7HEZmofgLaUAGn45
AuKW27Y/UCCJ4VHhr3nrqRMClCuE1lVcZ5xsqUlOqgYjIVZn8j9gXVJf9sW5n7PB
fTxF2S7I5HeEyu8r9cNkzLQREDzT2AUrSd6L2yCm6W/m7ZcTyoTRfFfB44S8hqEi
x1GXobkR2QqAqhd6gzIVie7JToM7FgXr+x9Tiv+ispi9SAIB9awHYzwZxm2Pxbz6
CMRVHZ879zlcxUc1ZSs+ozcJFsHLVYpscxdd7vUq5cDYQdHK6Be4wnCHIQIacXZI
AfKOvOwPWOJMONKzzxX6f0g3MVyE30eko6kkpq5BhujKQwWRTdlPwZ+eZUNW6BpM
qc0KxD9pO5iBN+JoFYUNrAqO+1VjuqG5yzj5uwkRijG0fzi6oxM911JQevuzweN/
DvtMx2BFYtL63N300CgiwhwRLxis5AtHjqTrthuFAV3zpTokKR7/YWJMIa1pmDy/
2+LKWAEFcJGd40g7FMoBCxl4s+w7IetHOrVQ24ve9Dnw3Y2kbYTM/OS/Yx4mZ0on
GQ96WgeAsRvOif889SFXTQ/fjZCL1ElRTXP2Cjsc9+BnmNDBm84K/tIozUNgd81P
taeobfhMOmO+X3Ikz6GaHxhaCFQit5jGIeJqXt0kvVUxkt+7du1+PasdMjiPPQCZ
Xg4rWoB241Hgwn32d3bTEx3i4aqUBSjuP5Gma/+0wS8y6Pgtyr3PyUC75TQC2j3j
nb3Xz9g4Rhk1gMyL88KGLRb543DENiDH1dcTee7Ke6GAhZjiU+YxDx7jhwjbY4Cn
hHhvicibNvbnV7c8/kVUvI+/5hGGnOx7S2lXDQKnpqOCJ/eAo0vfr7j3mCar9v4C
Dl3l588Zm/9iXmxH0zICBkv5YXLH0CnWNYG+9S18gnJLbYcdlJmstkSmjFlrbJXH
lNvXcty9B9+1E22Z/RzLdO40ZEYOpek7HBTYUxy7cSwpUV5twLuYAhtpozPTiJ2G
OipAD9vXfZlgR7ZjLp61iBftM06PQlmOdOLDrNZaw4zSpu3SwAhTkCzrsi25y8Fl
+Q+AnMslmsRPtcw0sek+oO2BIkObqXsvjFm18gZLlessunBelanPYROKVno3wWuJ
0os7QW6wE88dNuHnflSwDTxLhYBzJ1MpN6Ed8dixlxym6o4BH9tt8j6KcmUXkGLi
u2N3EYyD4tOq4wjcZ01oGzCeZ/5Xht+ey01fHr159L/oWhvrch37t78Al9vB3Eu6
aKevExVurwyTQchb73NPxHnBRi4v/w8RV80lTUCt/MVLXDiTfZjRADCi9QAU2jDH
VsNwViMIzxsI4TGHTkIHnpUBZK9REOW2WuzJnL2afWnB9Qrkrr5nb0T7BEbKJ8nd
QPWKIIB1Led7k5lCQcaZ75a3pMQ5KW+1kJjU2SgEhnr1UT9WCqj2k7wZWnLTa7V+
vMLTaB/hdXO60URg/S1FQrDzmMiWsdgVeAOPbhp84mGLaNSSoFnUdvLQQea0sF7Z
vuyF62Y8PF6UhDUI4+5R0RUlEKA4yF+kRGJsHX6+ZTUs0l4N/RVrGFRyw3SF2QgQ
GHoEKecny6ISIilEl4vR66NRnJuQLyXP8qKHNr5KRBDVSPlcTrkRN1Uy8pfsOLia
dKlCXf/g10PDT//PNszwykdOdTfE8iaHfy/noO2V4LjskA4a3Sq7O7PvJL6lxJO4
/Pc0jtH9EXFd4IJ4api8Zw2OAD0MbNOQl5kudrWn3E+lSh2vw/sHy0HEzwmC5Ut4
WTghFbB1gOECU41F1be9O4Ov2kktaH75quTfgHiEy7tnBKqgDGxphzRLKNYd5N/5
cupNSO2hjU8gm3z+yI4BIq5ohpGCoi6Aeg9M5zk6Xz3mw9IkLKf+AM6ppSFXQxsm
HfVjkgyy3QHMxa9OLGau6KfZUyKdk4Pb6xsU/2nJmP2JlZjFhPnMBeCLCcWCeIsB
PZxmUALoe4HLsXeLaRzjISXQzW+HAVMBblUPGF33w1iu83mLc2wyEXRUSEzwLWeh
PvQOR2uLWDMVpSlqhs5udwNI3eucnMIMVwlvSIq0Qg8wgkq7JTh5N18Q8kbFcZpk
DMbHiiLbyvK1fTSrTPEsMpc4mGXabX2Bmq7CrMb2cuu2ryoo1IjVKnlvqFzlxKGI
9zg6JE0ssfEr4ndpytm4CaREtBZGipPR2rq7XdoLTc0MoLDM0wv+blGX50PKCiIP

//pragma protect end_data_block
//pragma protect digest_block
eaoppACQ62mQeIFLc0jx2ahchBQ=
//pragma protect end_digest_block
//pragma protect end_protected
