// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:54 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
PQYXgnSyqQWMWA8rT+08vtAbmgQiwE+y7OG0VubtWsFfViBA/3YV/h7eqO+xyKjn
dgIU7WAVvMTbloJLZHgm4jooKGqa5x7LHvxjLWODR+vGh8BTHCq2RHBuce0HwF1I
AcitZvQk/pEuVo5mh2mI0t9JGvQVn/VFnecd2IG+fWc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19904)
sPJbrBjom4Y3fyGKsYuSe8G2BiRc41/smo13H+sE+W+/liLY/ny+d72ZaQ0Xh0So
Rb8GtBirvZ3w+gWo+iPld3PQY+8yIZZjEu1aM1+MLK5i/yEG94J0h3MFcMCAflPs
r/6/gl6taX5zQhp5gpPM5ob1M/+PWvjkR5BbIcJ9X734BudOrPko03190bADzNyV
KlDRo/4AI3kHSpWRGuMSy5KtPLiz/3LPyhnhzV4IzObvD05UIbQc9xc7xp02mDl1
THEWfvJFKrDLwqoqwzRzR2+RTxwFvEyTWm5MyFbAEwE5tiOUTE7rzP3Jvg2N4ew3
BjlK3+mSkcCqzmk3tTY5tbccltVl5fI8m8eTUYJCrH2z6D+/GXYneiviqOlCAF6o
GPv4TgwVNPdUNFSlWb4veP/HfRlj55tgCQK/irrIGWgHj19WW36dLOmtcDSRJUuc
9AAtB02e8dEUOJtnofDqqBxdofl0IBVNMFfriE350yfRT7X1BfQptwSZTi2jwJ/R
0HEPk80ruCr3xswrerMX+Tk/JBmicufqJTL4JQ3SW9KudsiOHpkliqP5nU+0UBRS
YygxUhxcoLZh2RwIuiBjb/G4TUG6n23BEfM7Mj/pf/Ij1haBE3EJNMAMOfK+yPdG
K9WHUTrL9LF/3Mnu2+wWfReE2QhWXnb+6/uleeQlOVmGPYbHJkNuM1ve5bkXBt18
W+zule1RB90W+qHqLN7imvIeX107p2FJV2lkmWuFDC1YjexKmF/B+10gb+LyGz5+
7qRUpQebvJeU+rLUMs7mS0y9WG3ntpTnYRYaIuexs9Qpcf46THaWqFwsN0NGwXr5
imQfNhFpd/7c3emBSPOJTKUUOpW/qKuEwxeCb3TPNxFbcS6kTZvq7TAxDXvuqAtD
pYv5heaWl2ow7BEXxEnMGkqe5UHuaqcXV3oVnDrGCeZN/0v+LNH6sBg8oRnF5FYK
c/AH4EOA8JVlxYlSXzaTFGy/NWXWUNJDqVYf8KPKDlW3itDTFu12xbwgB2CNJHLm
1t9m68gRH3ZD6UQ0mdXjLFClkQtMMEF3gRi6g2M980lYx8OpfZuVcI7CE+XJBclR
YjB55LDT8VLRKSRZi/YVu1JE7MCXQoYzC/z/T9UtaadC+w6TNFKEnSzHKBZrQeF/
6GyHqaFrTzsTtByX1vhMhuNyCng43kLGCN4B7vEjKxfo+xNiIpZcTUaY26PR9OmO
NyGjJRXk38vPbSp5KPNwpX99d2zZHdCEp5uYVWweumwvL2Sf+6Le4fqzP4ESoAkh
Yvoq9wUl4sN1V0wWJIsLvpa3NwzSXr+NMqem5HcGNsJZDeSlUaGyG3Obtfjs1eEl
xWkQ4zWu4N0Z1xvqIKG6r3QVftbroWmyB1kc9z1pUTpshkMOYOU/fZAG8p/t6Nsz
eWMRIO/6sxqhgNtUjlLjHQUL8dDKeVtpCVbIoBtudzWD50glVLH+ZtiYlTp5OF39
wid/UiLXft5cgWU1oGqiOFgkTU0bScQmcgCXFxgDEOsdbBmKIY7cEUzQwVPpmK5H
xvrDQz5UcB4Se7Ru6qakz+GCHw2Rc57bMF4usCz0kohNadrnCawRQIcsmBEk465S
aqHhLE9SVy7BBUO+6X4hXsRWzdqZujf4Avu9NJi9rI1QR7GrR7rPPb6/wlGz7qCt
WiVqkXU25bX3AHgWhGbl+d+MOBGKB+aw58Xx0707NBEsPtx93T1/WSdwQnbrTDT0
Q2X+mPxlAggQe7ulY//HBMsrdk3k2FroXuChBlkIj7svDax69YmNPXOlls8hfiwU
9gpEA/leE5gOif99doGEF8ZF/goOzvRvVI9a+7m5Rdag+nZ0pfWLeWUAAnSDrd1o
IW8M9QP9RkD836YVoTrHitiNl1i1OOGKkVP6lCNIpB+/C5P74L1I5hgz65ZQ9D6L
gEBxPpoO/iXm9u4uJUC8Qk9p0n92whqEXzX0ic8e5MQi2+tMH7yhe/4lMaSCU7B7
Ri1Xihzu84+pkjgXP6MALVHmE+mn2fbqt40AmcgOeqTjhoGk90BctLlUKZAHanx7
ExmbdrRoqqf5HZZmP3EpYqCLYtCNwOfTBmbfp5aC50Na7FbZAQula3I/VCR9PEQN
0l2K1OsoW2cwVx1UW3f0Sp28UPGBcZtwYbCOv4uAHwHIa7sTAMfov+ox9+r5F1xB
eP+H3hXdkscwLQuVC5WuDQgpoBiPASGpHTp5rBmGACEMV0ArBE2FXqu4prre595e
wtEMZs1026VdiFVYamMybStGupbU39lCIHDd5OPQS7ugkMO4u5bNOgXTbtFqgQAq
HdRQhKOwEAT9QkIXB0sPRfHPTaP5bWvJN5G8uNaNd6phwxtepPPrzlsuYy0lCPKF
f3p1V80Szf6QvtnWRTg53vJqkQXCnK9AJKq6m1wER8PTmJHkv8QMKAWRdGZkcF8Y
RcUUGlgp41oz/DaXXhYRlvbGeM6yDnMSzcnEFTuj7y6VZ3xqYzgfttJIJ4l1smfS
HK3us62zgCpQ2yOkVqLyPhjPBkm8Hi9ZtYJVcx9LktYkpTOq4Ev0hvQ+a7BT9y8+
H3D4UPUZPacIi4j4Dj4ReGVgS/nYNR9NJpRfP9iFNuLxAADSSeWQgkJNgQhnpf/q
h0OJyB1pKGaTqonFSKIE50VLDsFaGfEwrKfhW+nH6JOO/u0qmqj8TIZGT27ww/bt
DFNkCOrGbI/wgeQVvo57Mf4s5ld1jj2jGUKhJF941TdYBGF/tRw6bDwe4ZloQI8l
cZ3Akj9YzeiigUW2j2G2g+SKXbgelyi9V2p0ys+NdRetGe436L/IvTeIQmlaosE3
uASE/dpTQDiioHoxEguEQgJMzjL75XdKcfMWxbeULIbbO5GxJZYID82xErHTThem
fyLZYuCs30TZAULUMBfLuLiilhWygx8z2ebNO6AePqhsbYAUpctXmEMTahS2x8Er
UfBjfHt58gMr0GdaF/7MMM9rUbkqRNl4OpG/xjNbbHVIK8S+smC6FcsVHoAHl0V+
2/Letdlq8SbA2dJepbhen7iu6JRR4dOvZ+ouht0wL8dcmqnfYQgYHDMNdWB9XTUF
zITgDzVSRf+t+9lBTFrL7skwFQSRNvI0VCiL8XbFyITe6iJbc0Z0arpxZlWN2MDx
m/qBE3HeOrNebHaGHXk30ZbBT1LGMNzaOSwc1LwTbo2eakxljy1qp8bFyTJv9v5A
Mu/Dgskz9P1Gz60VyJ5yhE93POqwxte/QHb5hMyZ0sXTF6K+otTNUGpBsifqcQ/e
C+I8eZKujigOiB9DZelYbbbEtGjnFZ0y2a8Xp1hDru8sLxzfN9u+63YwWnpV22sS
fKDUcUJbIY+qzFZFHlpteYDWoe+BSyYvxr7xjMz+yjQmwUh/AusXOKmDHc+xZoTM
cDYJ7bKPbSVlMCFA+TyTTCy65bxRJAyphvSIgBj/ZoIvsjWN2I35CRTkL4ZRw5UD
2mangKiQhIHsjd99kg1lWFX4QQhepAkmfm9kSzkxJXzeuXeCb/ihrjRW3xcs5fzy
1cywDd12J9apbfeymxCPgsKnsIjMWbViOlcuDrBTek3bbrd681FTVo06921Mror/
9xScFjrkBuCgb7tewwr033XMTbGHwRHidfzRuS9GJMQ4XP5lKb8vJ8chQyBCLbWJ
l7spkPExvNCi4Ht8Ktk2mC5yR5tOpixr8cGWsBjLY/5qNXu3no6HS5X7fbDghdgP
NhMx8lVCxXsPsHXRnX/JOS5pQV+QsH1XCexQZm0uPH4FDnHocVgqHWG7FwqJHSbe
aD9XyO8ddp5N+Eg7JMB/Qtb+1pHK9wyBl6MjZlSXHhohcsAWpHoTR5EfJHwEFhIg
YYm+EPu9EblxSeg/cQZNeAa5Q2vRFgRaGTRNrv6hV8rYS+cM1LY4N2fCqqYFM6qm
I8aqHglLgubMTdYtAV/uUjmUnLck3vdAvLTsKS63YqsBRbEr+dWsD6v0cOq7HKOR
RY6a1AilKZx36HpJfmL1pcPzDGcLNsaa16Eu4irtxfo1864o+3g6ypfm5X/TR+XG
zIAba9OMlVtlbbG9el9taY6nC1j9v9C1hP+wmF62Byhg3XREKHDMK8O9IDIRXbSn
/1vrXRW23zYo1L3fJb7O0+socyX00B7aqDtGjLs8gmxniVLDBHtD+y4GVya6sEa6
eHkFw/7xAEEc+rrRBpUVVVwV+R2f2up1ZNIgGHkvRWDg1xb4vnbwXvWWGkCosOZ7
gP+FIeLA1o4ewoUsQrgSF9EbJdlOSO5s+O40UsTvs4vEjw5z3lKyZFRz0ghTARHW
2euF/x7SaoTssJ96vsYqC8mtfKG5MAb5xvSqNr8rHS5R43iWID4I3OcBjSg+tadu
tUghuXl289+u927dp9zv7fh1BiqAN+GCfvBj6pLRQfRATPZpXTuexBJDGWuF/7Lh
+IA7Jiwe6+G0y+/MNF7qKBW9pxmGmkpZDT4eHKfacTqucvqAEEDVKoz1P4WGCiRv
OKuvNIo0rVlFEBAftRhpRIw2kTeI9KTF1xIaJV4+Xqf63bEfQq2HgKm2LbIYXUeJ
KgZibXZc+/nKEZ7q/wkegDwPFK6Mh40nQR4Vw6rLgpC97FlF2g1NMgUWsV5tEdw5
SFo+FcUJ3XjEwBoQbHkclOIboVUdLldtBLsKaiXsGUtzUHNyIWj0uUu3xZ5mLsnM
vjJ9Sh6qrHKy7g7LVaZVcvhmxKTfeXWCqLjE4NEpgqBDGVsRU3T9mxMRDAe82AzL
aqYRhoTQooE6SAv7/lFKFub2p2uUj0sMWohCr4Ep5jH3jCemfO1K2HtmvHcspyvq
ctl29VrshrAVe2ZplzhfE1CFF+NdL4+JKwMTpWi3HJ+KHepVa49NPNojyiLTfd2b
CFcvTpCeAGHYQDO7X3Nyy/LAGkwXs1oKAphiJNksqs06FLIgpdCtmyEw6Lxx/YxS
tMkEXPG3zh1xfKIANpZZZekG2pCrDragbfn/C/bl0kOc7m66FCOBrnovX8TWu5kY
1Ch4/JpE0okn2GTOypZofYAgS+VPwNYW8NfSGbuWDYRJ7xcaEncK+TkAsZ5beFGc
XKj5FskOnv+asxgrsjCucnsFyudjZG2C72jVLtRjmOnbNlH9VZq1flhFQuccI8MD
Skn55Qy3RFN/ZuXRM5vukAqlS3yh/pgPWQz3QbFDO91uygutIRwim1QDXR1J49CM
eZVsKlheDUGKgedX3ZG3fjmSV1lngFLhHJc9NRdjH8e1vrnRiVl0k3GYMuEyihoN
s7rBVhUxK3U5jAj3kefH4FkhCR2/8JlU3dyH7fjHWqQtIZUlNK65CcyL+FnX0gWF
B/wANXjGlhFM6ICXUx4yVklKux9H5bFkSQs9YJIE0X8/JIsAZbpJK9LTXAWW0uXe
EFkiEXecrpeL17E/dqdDiddAkn7hIHxrrza2YRHTWoCn0t/D4rjv6n8UzEv2ywfh
0fFEOMHWFplDZjBl38nSQxd22MD/ddPglonYoZuJdiEi8QbWKNolhgwqJEQtnzuM
90rZ3ddIX7tKruOqWUtyHsHg++jDRa0vOY/xILZkYOyOz3gjxl67O5hJV4ZBd9GX
Jj8+xr8diUgvqVBte8ogS+p9eHrVzH7UaUWWjJZ/+9gJtekufSpJO0I5VdAF8fPv
LECiAdWe1n0du3MWN0n/zQD2kIPXV8AUPvJRPfaaOQDII3HmX+q5JiMZDXiKjlkn
MKSdFYiyGpu3/Kps6uT5Vk226NRstUAxHvMe40DWDr7+bXO2DuWF6LHgKCuj3UD7
pMv0tod14YLen7hbRmvHMNoEEKBReLRE6dxmlyyMONkvQONhl1dUe+oDLntPo30O
GJbdZVxhnf70Mcsa/iRwjNSyEYNJ4EJgHkU/GlHD7RHyZCXylt/XRyyT8lIaLd2k
MH6NjxmKO1keHB8EaJDJJGF++o5isEHG+VUjyiHlVfrE5YFnjFdSUPknFlEW10Wc
NsB+dcb3wM/cLp443N6Ux7goUnDTA1Pxz2iWge/+nW+SzzITWf5ILYgTFwvKxaym
LJw89eiKMv/JIbqXDa/HZtU5zpRhIhFuwjCu2xHm6GN713pr9ZfnwI7mLJRUNHBe
RgF5GJVH5zW6TyuRr4hk6OF+A8OAzkN0x50NBgBEur4mOb0c+1zs+iFuZZrEfzbo
tStW+x14UaioHMO1vCQyAZI0NWD6dnn8BshjxLLoGS1yTm7YKCRHwVmJrm+EmjkB
JC/thmLl/lvfk7MGXSIEUmvtLIm8S44J3GI7jpJqAoCHUIsJJ860G1RqkC2EAH94
++pbEQUeL5CjA09Mc3fEKG/D9PN95JM2XInbAVH067I5rJyIt8GHNDv/yF7DWnXI
hYU9ejTiA0XlcFVxh635J6l/sU4iBfBDQntSdlhPZJgPsZMlcix32CHBG7b3JOYy
AIc25H8c9Vi6UJu2MVPIrhwo70A0yKtk0rGxFo0Umg9HISOIMTpGbIyyoASMlb0r
m1Qrl1o6mYz3kVqLUqgyOYVDJB+IWSyWVhTgabVwRPynq9N/pphRLwTOmLIST1G2
LUW1O7AYU00MTJrScBni4Bcn46Bpp8Pdksmzc0NomfLiY8TH/+aJywXUZI6wVt1L
OhiV3XVI8fEbv1ozFr1kkL3CyG6UAS7VwDkLKhzaW9xaEA/0SqFk5Xyu0KxxqU6U
hcOVrQUnxJmhY05rAwjsGDVFDlKOQYwKt/J5FAQ+jXC03/o23Xwlk1Orw5ym5zeu
MCy31ztaobVuEzJ+GGkfthqfMpxYqkVRO5M8fjjwDLJ/EV3pwMp1UUg6LlCdgjzV
JjLypT6xn0npScXkNtgo2c8wi4LII73ax6rh7A4u/PRXo69qQmRSLAxTCixQVIBf
j3SvUf34UhJft+MfkCbdMMeWnVK594yeUTI9tP3U5rOi7EELdzlGbp26XMaNzl85
6jzf210mNilpW2KEW/yL0eZPv6zFmfq/E3wY0nyFtQ+T6qiALC5/ccaCaxpCO4BG
T7DIgJrNShMgqiJEeUNrbCVW9EHXYzGNvyq01kh+udtZgIXnxNZpCtWf8+HXbeBm
XIYPnuRq6QIYJZoi+82yIHHYsCQ1C3kAhqYWUcJMMzWLZ9VPK8aROuTF1ifJk38h
Mdv9bfXD9cZDbIworfrE0iyJ8HSWDn20J3jnh8Zd/JXdPN8Hj3pNGAUPQ90CfMJQ
njHGvMtY+xSVFl9VCIDex3N6HsGZrMwZOX97Rz2ksqjB3As6qJAkDJHEtVvi0xw8
4Q/JVaftyMUsX8fKJ4/s+kcp4UiyfUAZ4OewN/x2TgIVMua42gqd3HhfVKMT5Umz
btTFq9zSxnBLZEX3d8w1SLgKighKw9wja9rnX3V+FoIq2bt4K0HexR1C4RDa3wC2
m/PzaCKQzPvJTGcl5XwEvGBIYTAn1WeNeRpu2B44X14aRV27aW46FMzR9V+l0sBM
ngVYJdmSx4AFORopEmAF4Wm/tpQlXsw/bMLhkSB9+22ljGXefVqA4ZY0F+nEKYbW
CpM+01TM+wZI+fkNDKSVnFWUC+J4q3JSn3opnLoqUEA5EHdez9TtjZvIBdVMsV1z
gbodIFUgJuclrR54d3M5/51gVPIdKHrjvC7VEkRD6D8ZuQsgaIaE1F8JBzOizC7m
0hHn0K9JBc5O7bv3DM+dHvyfi0Rh3pBT05ziAIcT2w4cIui8IdyfXQa8gBLJ1xqJ
1XFOKn1ovhpQ1NZvePVDKY5X+NOwidXCO0oSOreT/XraSvErIOE6zyj6+0RVsOhx
MwJqgaYnOjl5Ko2S5zUExmngNmGFH4Z/Ql00/6NYgpzK/mUwhkxoPDteiWq+uFNU
9RmvACLOMaamtlXEPJWxTCVyigHN3UzKlBjRvk3XS6tmSv0F2t18NHxLqa1aHMbg
uSd1COQU3Fl+A+l2bic4Qb1RAJ2FEbdUb+l/OoQ1tiX/DGKaF5RHZSuNiwZKBA56
sQAInAoCQ88C9M44FdScPAuHIu4+oiQAN8sk1hSu90qBh4ZqyJJK5JvCCoUkWlsG
TyqukAhiICWFou11CIuaQ2HrvB46QG7tcHbUUioXMKprat/80PBBE0YDAoXguvS8
pQ6EVbrC+B02NgglyKB6cfhHGlNGaBB/68rumD3zdViiE/2hHaTgntCqyEW6TJ2r
lmX5I5pTIvkTKgwsWkQbkZEpq7fGnAiY/O/ypUvpkJPxThByC92JW676v3RLOzOf
rDX4p4uobRron5wWO15kzFedZ03c0ZsfS5hUuHSiXZMs/K9DtRw4M10PmhfU9YxZ
W9e+BK+riyrKasc+TdkawnZnSvXUlFl0VwqHBFQ5l2/zzZb2wRrPy3/gdeFeqpHx
REglIhGhds1EYp5ziD3xvpUq5cXTsgXlGV+5BYDJKuijVQzj8vmpimU0yHbmqu1E
gQbuzx+g+RLF1PMX5gHQnat9Yu2px/i3Q/cxGyjLYbt99G0LXtroro4shKBjSSV2
KvvNP/H9Qqoo0cafdMZCkgspwtr36LXxcjlwcxxmPQRvsShZZJyrB4D3oC4pyqah
z3nYx1GDmQp/zPVOL+djN+kLnGnQgw9/CnrcjN4cbVOww27Ctbx9Wiej21x0NDn9
lIQr3x3vamLV3VW1ttP+hXb2+b38jkVarSiu2tNwefpq/c6aHjwn5FYN9hgskqPz
huOoemCgLxvNkvTh1JbYvx4cmaBLUeSjlTySH9TWSCgw6CvDq4zq86Hyi7ZZWzRx
5SsqymBIQjyAY0cQJDDcxJYRocWDmH+YRlpspU+XoVF2Hp455ySTTUjPTd/G2H87
Mja/p1+rlWX4/UT0VjSppjFgW1JmjyVETqHernqI4dSsJRyaGJ9++GKDlAm+RE06
x9BaNKFvvdZ7ntxuHDIWj9q3pidwW9dqimddqjMG3oXK8HtIyOOD7S4UoUG2OUYo
63Rgi0HVEy0rhOILma4K0rlHeW6bBYvGVXvoSbpdftucCOxnBnbHBErtjMUgVwUu
aXYxFHUm+WB20/TgXFuLYDsyplFBh6oAi0ijLcmHKVDNiEuiyxQARk1GYL35IuVd
S9MFykhQ/XRbVY0rUOLpYzHV8181v3I5AwhhC0ao4yvcHa5N+B3mVqzWG+OxRSps
Y6O1jtkab2abruAYWBBM8Ens0FzZI7MAbu3h8ktP4m8+O/xxtYHmHp53X7RzYHZi
EJTgDae7vnNpo1BlRvJLXrbJPghj+fx99UlLafRbCj75AvX0+CLI+HReuZBAFHzI
5fW3n837H/+A5zvRaqDcI51H3FAlzbQiS5EL7T5BUT3p4f5VPUYJPWKo0iUW9vUD
jw6r5VQQHhxmrmwrpNKAGGXwtbXepFBX6dP1GvvpI673qXt2wydZvz2r7QX/i/nL
vPxKNxUfWGQIldPAM8oRnyJJW2MZZko9qYNv5LniSe1z1azyg3LZnSuVLsfoJukb
LBfebmpC22nyrawTRfw8YM+tVZrTFND7rmm6V2BpknDzS8rSkfIK8wJxQGHxFY0R
lIyzmUsZxzWD0eAyug761OY/cl+cMSGQMKwmLwNIf5RvGMa43PxljgHoJqMdRCnv
0qBn4zoKIsbj+VsoD0vN/CRhkWN9lkWgifboSdyy62MIRNZ9+IOOG4/bA3zsWB3p
UbahoFdewhn5/KqgGQX5GVd6pSz2kYXW5KoX0O1BGFCU5Qy2o9c8Db1xZilg9bL8
2N8c8rND/QKXdSCnGdlyDIVz0rKWGymA60Vzey/pueqLH+Va8W8x0BPkCTGgDDjp
bTl48ep1sWD6v+YHki4eOFfqHEinY7VWL6ExRV9raFukpdX20auVx8n0dHKbONF3
uS8chfHl/0dbV6yqUQgTtQnBsyRGlKWQyHJFqdExyyNzwydOE47eDUNPsoHgaJOG
O6WrjbVbuQ3axk2t6e0HDNeuxuJtDE93iOceX5AO2NK/38E0CjZMsL9yU3+0cGoV
Y+9ClJWZMJ4NiaTv47gXgYcnSZcJUVqur7TVD0QTysl01S3M+ZtIRcSbUnavA3Pq
OXhcuk2mxKJ4PVy9km9agIOdhT3t0XA8YJcGv3/Aa5x3D3KA0/wSZNLb8WSt+ElU
sB15NhXmw5hhLVyufuhjPHVtf4CuV2ZTgvlehc6FA25ptcWfMQjhIQwmCy9ERP1A
myvz3/2BmbkBbC2c2pBvj5F8AHRFKV98nIaiC8lMR7J+HB8ZRhvCFyZKeRMaY9ET
SFKyvj2yZxmdZVV8WQiVTfIJMqMbYw1chNYFbQjxcEXSVt7kZEbPJhU8wawFRJUE
F4uve+erPcmGQAdaaOEHSl5YZ0269JwLJxnFMQHDi//bMxeo0pKhQectkfSpaCL2
eG5Wg7qG9mcVsMAcHKwCeZgvtabk8JqhWVAiz33JFxQK8l2Ymjgzarkb+aekiI9l
U4Pc+zWODnng0oHmmpSdqNMLLMys74BNjCWTAX/y1ujbd7i9HhUrT+hTQc0h1ey7
/3NTsQqF7Zr7BYPNNf+P7xGr3W0Y30bsbOS0iA9X89nRoCpVKvm85HAC6nVUWg/Y
mIbSQmwQOnF20IAgIJ0eQthH6y93C97O1BAuvQEsMc5CIHwxE3uk5LGliYAzx8lq
EGAVVzJPiQd6buZd0r91N/Tvp3VxXFHqTpQha03VCbNnmr3al/YS/dq2zr37Ojfz
hsVHofQs0D0fhW6SCBCIIn02gxyAwGyIW9du21eBAUWbw9hCZgeW+FV3+EKSgIqh
/TEGY8zI2r2cjf8Y39Qh+khmct8zS0WBxWpTrF60DmYmVbab72ND+FQDUfOjLyNj
iwFNt7WF9sBvX28gh9ZmtdXlRzf8fuGR4CpcGaOP5MQEDqjmJlu+b3KxGm5gCwxa
t9cKZWSFIh2eIHJEfnP352G28g/C/cUXEiPtX6hz1GV7n0b+VfQTnxYkzraguKTF
Vcm8AQRSRojgo2QSJ7Vj6OsH8dKIxfHSvnEEHrUrWapr3kmU+kni4fkUc/EgBTiD
2IzqaXVonV945oJHm5FXcknYqTAIvzS0VDEhKtbiO/01UC8sdb3wwFC7bsFHY6IV
AkbTipXGK1a1jOW1vmxXABzLkgm80gjyhTVqbptQuYEDWrHCSbSzI+uN2zRjvEJG
017dw71Px/AfScfnC6iHZwUNdWk7UnmJEhQeGUFnVGIzBM/6tgWhjitlK/9LIk6U
ejdLq0MNrXXD/czdcmQ7L115HByo2v5T3o57HnZpN9x2+joFSL+kN4VxzbHPBJQf
j4ox/b7COP2ZpoZbJQgOojYoncnQosK4q5yqm+hiSGht7f0qv3xzURLn72wyz/T3
jd4po6t2BkbOrzeYNGV4i1NnjZi1pX2h97MpZRehNh5ESySoGTQvD/jNFH2aPJws
1wOLPNqYLYr5BVByVuSALVzVIHS8hnkW+kjVDuFtqIDvC2dKU7p0hJb5ifUl1lTx
nffoS8cK0AuHLIwR+Guws+3MCRSC6symHkfoVSHtMKcyasa3e9RNoC4+2jyIZ+Ov
xAAyrDZOsyLKn0LUb/WUXOIRqW1aOZ/oc5I24k5ETeJCw7Q040dXCgmSgqtFQicv
ZIJvJMSJuCd4aAIznuIXlmV+FOHSI75p+J3Ftha4MdRExzEwp6jsZ41LILo/3TvT
79ugO3v3CX9+oydLSbF+QYA7ZbMJtLSIarGXUPPZtJs8XQMddrwNmdISdCaBXcpO
CDXi7qmtY2Nj/s69jGUrejQMAU/cm5yGvE69cwtCHSQQDHVKqgZGHcRklG4wDK99
d588W+TEnXZmwUlwtdwaGs7VVEyjhCDeIMXmczY6dlX9T1vWqE9F/7xyWdfHHez7
7AgUsz2+EVeXnK/xyEH+0j6woKm9QmT/5prPH1Ut5Tqe+zaBprJJsta6ekTQS2T2
Og8CcN0PZnOWsDyOgfSqDzWNBiWpkhpcZAIrVEVtG347wvsz5G6QD8C7QWXj1YI6
Vr01r+QEdp4tfRcKw4tIgqaWje7qHPCtMErtxmfHpm0jL1LuKhosLR4jWOaXUsxK
z2qjLlI3g+ySJWXsbwV8A7/xhpwJNolPIOt4LlnVPrZ73LwXzWjzU5w13utHn4LE
5GAJY1VPVsLfVnBpHHQ2lcuUc4S0pxpoh4vFk894Y6p5TxR97gGOLHi6puhkiIKb
p3ClIU22192loE0QHChE7Q135IbfTi4AlAaMOpqt52t1JoGW1f+Uo2hzs/FHeW/K
s63LqxKFDISLhbNCWatNyr/u3+xBKtNOt7FCpUxCM/xlZFgd974ntXImvbrHBTTC
RDmMIIvKYaUArGSY5C0LC34zqPLp6+Gm1yrl4tHSe1kCpPATCwQY9LJbhrLpeyCC
mZJBSzlHPxU51LSWBDx1TbD8rmqJ/1vhZVW3VNnia1zxkSTjQY9/8X+Z26qPICc2
3jWCH2jpHBGPo0HHXQRKIUVZwtm0q2TpDM1n4kX/qOLthKjDL6aFGzMoUc4OgTSp
aVWOFGsprHTrc7Tc4UmjFzrtJ30eIwDHRESDpf/2gXpqa3Doc60lND9GB5U0oERK
/TYwiaYTETzfimWe5T17wPERi4EYtQ6jtBNT5nU1/s3ePLK43tVspaillCvC3xYg
QJESyr7Nn8Zu5UAJ8NWu4vuSUsLMfwJI6Nl85g0sL6z9iaKYswECpKUY98b9LYn4
0blvW7kzNmYwzpRki2DCSH+SV3qDUgCTk4jzAyjQdeZfZcG6soW4hAFwYPhfViKO
XFdC7V4SJ2Gw3ytN4YFmoB7vd1jrp7r99b7P905Mg+y3EFE0V+Hc7TJa5XOsethv
9xKX7nHzXd/IIiQhHk/9DZ1sKcq0J5nJe2+KTt5m7MUi/rgQZsvev4CAR92TgyKa
9JPu53s3Renhu64xuvecxJF5NTxnyFJp915RCP4RuYwAsFUyGTHKNGUDKO4hIeCq
09Bzucxz7HHSIyWEBzOB6ubYyU1MiAF2kxC7RexsOQbZYt+dxcWeNkWObF6QRCRq
orIoL3ZNsSWtv4V4tHUWhFXOypAWkf2sxQt5hw6jcrFVg6fhDq7pe/5HRG5ayXaX
PjxzgPi9ptsC5BuJqJvkAOJuC8igY1Zy5g6NwL6pbmXJNpzeVWnJQI6hgaOG4RCq
v7k/nYE/sYojbdwjMZGZA3VfLQVZZJcYPmgUqly3ZGgQeJQdS3ZmhrMs9cn+t8iH
ixAtwoc8EiYBL9VoYFHC15cLlx+UC77+Qi+npoEr7hqT4CNEx958B/MU8sGGO+8Z
Kj07vnDtFNaDS8eQforsL7nTuQv36aV8NGEhegH4460fcQDsoW0tK+ruL8LkwFBI
z8SmD1bXeL/jRLMIqDemR/nJNGNz0GmByRB1SL1l4fGky5oIK79JVRL9Ke4GRfIL
8UobE+6/59G2aYzsOGnmAGD5Qtbj234eTgZVvGScii6p/NCKwpiTdwkZIjuWJc9Z
oTvuY/NGXei4gVy7BWp4JlOgDecPweY8NumK8IpQOT7Std4R3qyS0qsa8mn03Boz
qYy256AU/ihpk0C36Z44nAGcgPxpkYWhryK7RSS8G33ETFEW/xjj20t2iJ8MEhfW
I4Dhv7CPuxKO4fo0tTtpAbYkRVOqLBUSnjTixATAY1l0NdkGh1U97j5xPj4JDjpV
SUIbJ2yYFXQBxG4DFE6Ot2OXM7jlBHwbsVBpNAgwtCy34FQQhp76IgC4hkXJ55/v
UN60eIUZP0KCIXKwE7M6lwPUt79gYRXFs11iCeqZfUISJvgdtfGap/j3X9I1yPx5
O18Ai5++u70D7hlO7qE4RW2JMLn3gIR0DUWOX61y/oU2ke7lpqke6iMjq7C7HEY/
dYX5jXrsxzFYxhLnvK51wD0f/F9+lEPBX8ANqQPrjkr7TL+TX/1BBNhVs07AYWSE
7Sg5GZv4oCxJJOlEMiAnViV8UtR5w43wXbOHfSrM2Kb7h1mnu8Nh1YwD/EtCZlqb
99mXqQNmJX69JQcGh3J7KnoKW9s0PCiG4utvNQx9Zx9hr7EI9CsOymNfNgQgRw5q
csSrxZXvVzknhBKxlfMxBIJLUMCfn0xa/th4kZaUsaEUTKxI69LKSYnCG90W0VKx
dXofDpp7iIOqKPZw/Ef849uVKwjufV3SpgdNZNAawgekzGkg8bPAecg2NvBlMO3T
g7F/nCLa4Ny1VshiWUy/RRHPvfh3buILdOZytRSKGIm6d6ROl4vOP4dxfKOBIuVz
i9goO993ljN1bJWMwaD4rZQrUevPv5RQzOx85P1lnA+qHEtOD3k+qyoggXhHt7BE
XjCezn7w40GJTs1rzc72XhiZZASnrp+P249PaQ9RInKuFD9jS/+6aH5JsWRX8SkG
KtpAUDVzV8+MwBZdMXh6ZCmqA6KACooCx0ddDpZTBrFW8EJC8usy6dd9FFrZt6M+
oyAyj8s25EWOvRbFulcXV76Kir0wortUy85AFTUtpCuzx0NssvvsXqWnHitp9lrl
Ams2P/Vtp2fV3wRMKu6m7IotAmcIpT9CSuWlHHopYkb5fOeXXUjExjo5WYsesKYv
EgFdHkA14dHHLaWvzv8msxGgi1cVQw/BPOGey/a1krczqo/0ilFiPKcUuCxHhyFS
P6wKEwtbmpA9YKBE/eEUlHHtsg3V7RJPjWWXZWUEgHGk1NtSpzeugbsGkM6aVG26
mQErFcbg7uzfbTtb+dGxmuoagek7T/7MsHi5OgJZ5heTlehTfp95rmuRfo5k0Gnj
HLAjD2yPvbVtQlrBCHMR+1bhNbUUin64Zl985lzLM4/ozm/3mWA2caC0GJxJ7xTA
hNnWYriKgIJu88O9DzvyaW3rVQlupM2rQT/N0RLBuxxtDG06BmBKnVIZQNjK9/2A
Eo5elYsy1xjbp+aiToMqVW9W5aFA2LRPgkY4Hvlmle+asR/8rkevLxy6frBtD0zZ
JTm3Mr090B++mTpcUHsfhntCdIU6+VwklN2NcGfrLCEdzqScO0i1A0hkRQxyKQCE
k4xnMoI3c4hGUqIMjS0sQFHOScVFebseESfaSDVSU0oGetTJi+kwdldIwlbkqU7p
nSjgu2W0r/IomfX/Bb0gumLuW5WmOwnnX/kQBSI7zitQdnfDg2UQx7q+uRUZg1xm
Iv7BE9wTTlMTNPeCJn7qPyYI6zqcXJ0+AfiO3Y1uhfxJ/+hbLfH2XSiU4BwuZ65V
DdPdFP1QidT4baVY5mpxkix/atjjJaBuOARuaiRFGJuJjolE76RcvfhA3Qx3TUTO
sI5rQKjN/JtlPF19Sj7eD6BFF+ddr0iFYEzUkaLYE+hZybwgSXccLtJKt0vD3F0i
JfYlNLjD48+f+2PTMMcSvQ8pC4bwd05FtkuW9XetZ7XyzclHo0HAnq+8N/17X8lQ
Lbb7Q8lfDUByCMOe8DSqC+83VISpS2Ht2JRyhHMbZM3NQ0o29oLMWVNniMRTEi2c
8BBj2F7oxxvmsfwxyEN+M1uE1EDbbnm1vdf7tnE0S3atF5rWoKxq9OW1VD9INH4r
IpoNzZAXY47Mpa5JcpBVWFytCczoMh288RpRWDNuE3NwQBuzepWzZer4slf1E+P0
9vtNwCgnetgoWY8nZ83z43B9hWs4fiDk+NZy77Z/Gm2WzDBL2CUQl+F/4ySJYsBb
SWVXfZ992Psqa/zq7oz56Qj5DG9KhfNxiBFBsQjNaH3+bHSHA+DKtneKHv2A6IXG
cV0C6uqcW2w8DtviMOtgNqouoM5LZO+pfgDTdqC0eHgQiVdaywdHvrT1tJLSTnY0
TATx9qcNq7PmC2onxgy9Zs4VUTjwhYKKDcXO/4mGIA6SFoMNpnPBvG5T0g7ZxjjH
+SBS7PNPBZisWddoKwzu39VI+wryB5X06g6FWYy6Ed0WTi7WMs5oXcQ/UC7YP+Qy
IgMicVzhd8kIgpQzAFFCN8YbGiEcsqSpaq3nlGtUVXMFdEHeT0Myji86HkWoeqRc
CgbB2H7JRXb0D9+V2ypZeQryVXSnuWwptKn7VDHWHSWMgITZUQI+jhZIAWr6ccIY
9D7DDwrYFHUF6tD+Qhx3qidKZ4jg2CLuk8FrC2OrXSjb2mmouqXcNbUGHM8XAM9Y
ttXPG1IhwR9aVKpxnLQ36Q2CebTHVgeRzl/4qxQ2nciA7YoBW7f/TuDw//DpIAW7
ckyK9pnWEQ5+ATOdQKmGZ6z0Oydck5fvebdeAZq37x7sFprrAzhUUXoWYJ93HBlx
Yp46qlDH0jcVU7BfeKi7lnVJ28cju8b0DrNmT3PBmrLmQndfAkNh8TDX1q0UeclH
T96llxxEBcj7UxisoMgLNgrkZo01Y2BtRWNIen+1XW7jP/sf0xB09Wv1NRmJyrl5
vQkxSElOx+pCkJZMmWM2OEgh4OGsKm50VVLlxjAa9ZV17a4z8EVBkFZMKcA2vfT5
McuDGXiruFsYnJN9w2Panv+BN4+LJz6GCInRmE4HlQDCHzLjB8PlMnl2lLb+4tlL
BrB9BdSVA2YQMircOxPT9shC/kxvHamgVHLuZDja7mRsM4upGDL66Uk3Oehrp5e1
jikBEfspGlvwARc6wpEnT9+j40gsuCBA7HoyGGg/WGXir5eQhVdCTLVcW+JVxFOO
pWhdz5cidXY4+FOxRkW3wCjr1SK5N9AwVSfhQT8thNGqhfon7rQ93Jzo+Ir4Kcmm
MBPE051skqUXFfJGctLaW4a6+uINoOWbdWdqIY9fx4C3bIc0Py6aGkJgCMJgSK6v
W0emx4wuZwbswwMD3ViVH+HpFS3QcralkxXnfDYrO+dQ5ATITiPW7RaxWgaBcz5W
HYQSzTnEyqCglsX+EAWJXMlm2tU9vaJqWI+WBF+HhoLIE3ECaK4B3m2ltcPiY1sD
aF+DYYIy7a6NZIEbawUG2AEVAVlnTTrnGt/XHML+aZpQ1unS/pqaG56USEbjwD5I
ALfa8G/sb3cb6DrnbRSfrapgTzXwo7Y4Ph5DYjMatW3oGxYAajP1htXj21Dx0lOj
GfCYh6bf/tUqOpp9BMwDCRX4Kw6M5vmE2akZ/t7wsQTKUkpS1sY34zCs2/aZ/Dsm
QIrW6IRIpKuOPRl/wnoRCWjRV/LjoBMyYj2372lPgpEeEmN5c0REn0wRmXNKIR+n
uT74ozLipAqwY9MKAwrHcPfzzX5vA6ZbD9tbZGNzru7OVqvr8TnGKxzfgC2XwwAa
jp89QV3x+bo2UjtgvIj+ujjCZo7iRm1q0HHYdggwPVOTblupA9VtcIeEIMBQ/5RN
IbgZralFAfM8+hz7zZHG0ZJ1RH4ye0kmnA1O7OT/7daYylbwL+j6JzoVJW094go6
GLf+cW+R6Oo/EVSoKt3p/lHnUhnWvuJJBYfAsS4iSv3Fgxviq1iFwCM0Scr+9Cse
oxZOkJCR1BO5zAZY/nqVsBGhz9QItL+jZ58oxXsAKoVvpWOD0ZeNENNii0PF4g4C
W529/eboOj0VX92dkWqXRc02c4MYBdVAeBj4i9C6qNg4iRxI+0dUeTtCXrLzU6+4
F3d8wye0IPcjntUwrYfaQWo3yhRILACtpE3sNvDZCV24yHgetfsI4xmseOOtZyLf
i3rfn06FfwVJ2jAqVZtXcCIVKjIEg72ZOQCPOl7mHRMcL5L0ug2xKJlldh4V7me0
zRR4xetnM1dfNlvsWVyQiSsSXMR+iFVyOf7uQJ/bbmXz3JHljrMH9EkWBrQA6JEy
1YlZh+gsT4a8YYwF+fytKfnL0obDR+RQMGjJXemt/XhlOnGeusdzOyT/Tcj0BNlN
F+yveOdZHwheSRYIQN/6k7qfp4YjICnkFLEFjbMdG8x9gz72jmtNAdEnK42sHVr4
T0H4hd8daHWRZ2rA1GdNqdBD8wNE29NkxtQokENV4VtA0QNir5v6Mp5Hm+X+ifSr
vt0MeV1dlMH5C0el/AgUK2bub0tmOye1SGFc+AMHCnxtOD0wU/EG9eMD+3UheHsF
THBbQP3OEuzzjWcfwptY107ZzRLNI2ELu5b0KrXo0AqB3HCOM3HNasEgsCe49Pbz
Zd/RNtQvZV4rH0xjDdSV16nKAwjobRzzknduGcnTt+xruiOncWVmEdF91LKxNT+N
cgLgLfowLQiaetSZlE6zkrDS0FhXVT0YFzeJcQBfi93Gy3Z7hbubY/tw/py3xfta
xxdVEOTauoV8bLiYCvIMMCkrj+aGlK7cIGkEXZ8v3c2u523aWw6TA4uaygYEtJ/L
TqhnWHGTsztJP3Ah4INQjxBj/S86f4Ym1Oo0utnIGeL5nBduXwMHajASqSZEqa88
L6bxx9mAoeEoSk4rNlXf251mfaParoXSPuUNcQaQQihdOHv2hEcJqOKXfopFbLbj
LK5k7Po0xXt7jlXh0DYoPWGCraxC+biCJro+mgWyS6prMFg31mzafEHNqaIg6i7x
8BwX/gBV5cfnljlDoIEcDjOZ0Uyz3WZyaIUEnVm2CKqBf8zprG9dzdJGVWNgbXBZ
IXDEsxzyJLGhqVw/WSUh7ZEd5KKxx1xg57pEl0onUluB+e9rn/yzW0H4vR3mLGik
u1h1nXKguwCLti5C/E6fQeZ2yc/a/qNTMwt9htx+FPgx15porBlF5+tA7dWIL6jI
1r+9QQQnyF0oTI4CYHZKjm9ExbkP1vMOEGmZplydSXIzZk8aj6lqiX+pNunmwi9d
7KvVm4WONFJ8TTCESYJAdoARvC22ZYOCxJkdzP6CCZukPJyBoIA4rst48jyOVAxs
GfjZiALxUXDtnVrrKzM6UXqepbVpgpchNhIDT+h7IB8h1Kn7EYOkzKKPZeNC5eRz
0u/5sqcpP4PiD6aAmYRz5qAHILBqvWEZJh57WG4mQxCsOrxkkOnyiFzQDxPJEsTa
7XqPsA/JPnqDrioN6gBsrRiZcBbxihIb8IdKoMfoVdQuphuTkkcFu8jbKRuLmZG1
PtBdJKvtsXzk2UT++vCLG/pNoNcaxROVUxeAkW/0TJO6nevFgQ7TazMrTGmFDHbf
6i5xqodD3ua05J2NUD7E0Aya0DOEIgqjtt87bZebxnNBQn6BMCmMi8Y/2KonlwCm
MJRh7kczwaP4ZOUYEcMOJQxZKG937oRSBAcpMszpe+Mt5s7X+9IMlL9KWFLjvXUj
CkOjhGcrqRFVOlDjKZXs7kh2WEmLMMQ4/k/5AMc4BkP/9h5qoMXI9dGgG3XYLlz3
HhPjy+7TkBqWU09q8k0ZfOb3e7dW5hBXFODXNOF63wD5WsMFRB6NqC+fCQVFiv/6
XKBQy1AxlEDIhSMbdjnzHer2B4QDuGU0Y9xyIZQ6/LMdDM//bcZ6LQkV4abKhYtz
b8KYbvrhLB4pv0IxqlO5F87w/cvu1ua060HlfgttzHE1n7tXF0i1731dFwtWB0WJ
Ywjxjpyu5ak0ny1OdHz8HJsmNzjkEr+h8YfKKKRd0UUox+wtpUC4zlBrdUKLvv8l
tJBPSJAxIzMehQWjNqrJgXRkB2j9OLsZ5AQebRP0DtGQCCkWVPBtmqj2/Mq6p+mw
T95VyP4cUrsRZMzvvYILqPo1/qXeqWoiFNy7zwio5e2wWykBasB/efpujjaAt1iA
Ho4zeFZP17yF3IyZVZzyGVHBucPLBy6taYg2nfvXe50sIvPuHyp1AZzwgH9lhqtC
Slce3ssN66C8o+lgnfsPYZ3efekl2aSd1x1AvfnLKFWA4LQJ1uci/criP9PKzRbF
eW1ssp3cCrFu3YHHB2Gb3taTF8XjEQufPXLxABwXugk3Gh7ra+7jym9YKQ+yJBdr
6mAVrt4r6DRVuhhlluLfskJcveNWPdLtHvvHi95JXtg5R2llt8oKa+axPRiYuov+
g1ENUE3xxHcl9vMn1YKwfHdS1KDmhJi0mKLMW9N9vbmN2uOHpyKOTzua7325I9uV
vET+jaKWcFtexsLHDHG42xGs/hYUqVveOsgT9OVCqXttlwx0Z6vUiUcVyIVXareV
gBoTC5kDzPmxfGW2pcDlO5hM2RBzqltKK2qLjZ012SRTeERRtBoE8lajdy5l8GiR
k9vDrXY4Bv6GxWgQGcjJKtCkq3IrlFxNxpTuSrQGWL/rR165fFxXLBOZ0VJrAmuZ
Uveoo1T0h8rg42vvJWkRWkL/r8f8Bt0h7waRJnj3Q2ZjNTFlzfmUEs17LDhdpI3q
3wfGFgWOanfGme+M8OQ3PMx2fmQsQEHmA91av8NeaffY9DBSqVt9hjG6uEyGHCKo
HsECIsL3OlikK/J62fxjv2B5ZR9hhImm5HazzI3ATmdQ6ZxwwXVDYmw5ce7/k2j4
6wLufEsy9x97uR6KT4ajEoqG6ViZkeV6no7ueMT4XXJRZGI2iyTcjYI8qM+3S/MT
6F+IeWkQgWudN0HMGEUActUCJew+YnioMgMkkNIYxNvmUM4jSUwBwT5TjK1qxm0k
FrszKTxo5TELlDbO7UIMRNf/5jYFRW/XHTTycF4asKz63kw69mft0ggsHrHs9Dne
+GgXPaY+Kz6qrn7lRaIclc/A2wsHfuKaO5uWZ4dZRqMpI0IJtUiLmtRnRBzRgAh9
I/+tpPAT5g+g32p8vzhEmblx9XVkKskmfFmgJtFUzGxmIxM3EZ6tWwZ3LrVRnY7B
Xk5HqOmRmnSTCSxxrcjVTlKc9g1LbadLSZI+Krcnw5qCU3or8AvYstNIZuTiP89/
Fn5RS9avuhvwvssWWAg3XsP74+A666GTYxeCgPiRg8xmcO1nlN/Ex2V7idEQ8epN
PA7CXzu0HIDmzjcljfdnC0sB6vVyfgDBq7ZZ00lM2UJk0bp1oO36wMRlXcG1GWyq
YzMPQjfe4y8ikUb66yjfRvjsubzHbiyWORtkxLULZA6BxtM8qRWlw2rW8aNCG4e1
DpwxX90b+9cSNXdUm2BqzJjvJUtccjbbAirzYoKpaKNlgsGGKQ6SyTMo4piuC4m7
twVactTKwq2nyqHigPXZ8nOa9gi26tLfmbRYBYl2jS17mtzKrOxSwB13MyJ8E5JQ
yALtq9IAxc33eXsCIg85zkoNfKW5jeARr7IFbbGIMVxd/rzmY1exA574D1/5hcoY
fNQx89ZRkYIQwG4bbLAhVVLBxsmAjrZQ5ElDUak7NOhwfLnWi46yZ4lPRRDRc6CS
khEn5/BTc0MLrXGP1+J4OYTzHbvX9RdtDMrcP7a1fD1kNsJ4o94+0oLoRrtIiIeP
8bsB79Hsex35z8okFgxFKtjXoE6Z22UvTXNkLp11eYGexRXruiVCljF8DZsuRaw9
Jyx5RHwX82LpCP0nZe9NdiFuRhGR5kDjj21CzmQdfcp58b06umKg0/nmBqfq1AnM
YOHngq8zkyxV1LB07nTlNQHHDyJgK1DHbVi5MsJpqg7UnVQXk5UVGO+tuLTYvyb4
mDk/FCvjKDiFtXk/epOzGlqStz5k5rdx+bVng1pwpbWnG53S17ZzEBqKhlHOmcnl
KBvgaJCqGYhSYSSCPvRjsUaexz/tKcTF/o7MDR5vYULgrjJ6LglJPMltxDogwQ+s
F1oNtCH2IQhH298OA8+DIVDALeR2NXr2f51WlL1Kc/TOL8zel37QU0JrluX+Gwfi
MTXsoxL57TTWFc4xf/4sD21Gx88MLAjTunUBxQWjIP+sDFfNW0sclGPHL2eofTrz
yBvyFY+QaSCgvCavBJXzxJAGLKfNJO+jtf/VQkCvkEV/zPbQ4SNgczMH0DyTg5tM
2GyvPHWMDstw637o3Fpsjx5tKDA5uek1gA0zAFruXVxI7rtPwEoHkDQFbIodjtwP
yHoY/56Ke1C1y3+hdkMQdDmm0XN/fFpOQ0EmFWh1RCIQI6JpNB5XRjgFjSTE2S2U
8NUtnupFxEOGU7td5KIcCYp6y0lI1B0Ah0VcIGuZXxr6Qk0I+Gz2Fmt6oQ69yqHh
GC6SC3JW0YlApR+6YrZ3lQbuuU2dPuwccnHDFkYv47elY2Jbd/PwpihcDwTLzZtH
BRlIs+rNYpqUxMfGETVn3iy488QJmTJb1hVQiJ3UpwNC9sk4TPVsxzNJW55Urp+P
um1BblWya/o0qne1t7Dy0/3toEqFEF8WC+FNv182MkJUu8W2qnH8n/oOtBSY+tAr
P/NavInBnkQs2zn/Q+PRD0J78j8sdi3jgHN86pa9mlmpHgu5syDSoncjzzGytWFy
OPXfOvpm+xuf3r0X/tGf4zJuRefnMsv2iOtAGnwV9qYCgHo5INv1dzhCMbkG5Yf/
jd7NT+9aNfJGw/qpJ599+f1sxLdnS386QunbgUJLnNKX5gKIVZLsMdb86RAv20sG
iB98tYpmKL+Nt1UfGOAu2VGvYCi7bUHR/3DXp5UAD0NWk+1j302NSAuqBGpZ5x12
reQyRgtFQnDEWmQvkGp9AhX/g3FX7+VfYrBfHMbXlZ1xeVLJlw0qKrjGThN6bxeV
kNNWPtcbz+K0dSZiVwipdzeRag+As5Jm1tsPpnsuN2545wBh1IYPpceT708bKrAI
s/wcO+CgST2sbfGjj29Gu2yyHcDfxd6TyJENzD4M5xngB+L/xqj44hz6+D1HyIh3
MS7z4HF44fxp3mfTMCaWObRlc9MaEdiFQjasFotPg1ZwUUei8vNgSYxL+AevM1FJ
MJC1rXJUyAAHCdbdLW4HvBn3tEqDOkHb7xfmhDCQnk9r166v08IbrrSMscgn5S9+
dvNwSQG4GNbyybkjysvttueDasW1ACa8pTbNKMq7TY/9kdb38xadG5bkwhWku5pe
7bX3WTnvkcAr+f/6je+QzZRH2jTHA92GseJS0kNpiKUp/l1sUwLNuhj6B8zIzJlu
dTcpjrX3Qv6zP/oos2oo38JxPNRKT2Vod4VA5V9lOUkJaVD8NA8R3DvbXPSAuLyt
PYEwfE6hEEu7Wk+0j40hfW7N6QOk/D/jaN9glZ+FEM09b6nruFqRlFAPQ0M8kdJk
Lsv+Ny/Vn0p4PbAg3I0B/2eoxwuwL7nCADJQxi9+we6a7l+0gBvQJgPBSzfXFr97
T1ny0L3zzRXv7+GorH5T8LicgSTFEy0b0VdYeHP1Dy8e7Zp2wn02Ux+tfVhYCQvv
eRft0lkknUe0s686FQzOZ57OR+0nM8wIAfEMhcBUwxOl3ehTQKO05CpMAQGIWx3v
LBYyOcGXF5PUcNGoc5tMYecf/2eDxBD2UQjW1VJDAnsWDFLdKlevcf6SfX+hmmSr
B6VhzzdEnBQLsPmTRSuK9UaJIMmcGMRNfkTAZWh+JOs4uUV5qHyxkNPsyPSvRZNo
EMXeaI9AjdzDUqGBmwrPxFHUTFktDemp3/nvcrNh+r+zxiJ+/4M9vNFf+DI+0NBA
oud0ZX1HwcJjtUpu7leRGTqfA8W3acYa2Lte9fMAKiIJhGgyGRArzNdHgVBjaRld
wKaQW6UL6S/Ypt1yNeRlL3UvpiJ/IJkbi3noTthv64yRIe1TT1bSN9GdBczgaKFD
P11uHJHFWMC6Dz0HNbbc7mqLGNINg6UwB/1JMo0mDL3m8wOncNk+XU5IJwjWpY41
S9vKDWC6OI6xDURFH3AzaEjphUk6WdFNtHEN0dQ6wUXdQ/xEgQjyWtJDRV6iQ/YD
KQL9J3B/z3RUN0VE+l05DdrKpmKlry4/HtNgrceiasEW4m82RaL6r+bnNnqTLLxM
TPmwFOkrMASVnAj+BPTKefhzCKiLDE71xU+ZQ9nkneS5jh1pD/JaqepsVkFwsDpw
SOopwyy8JFx4YmqTq2QFP809x3wiJRow8Om2fQWuGSXNZTyzfPWBCeb7G0P6CqHO
khLuSjUGaPT2CcZ5qx1ZV/4zoj7Q1DKq2Iv4DCZBUp0pNJRY45THTNj3cMWsMeKy
mWeLoCAqTIJfNDPP91Uq7gQx0KdG5wIDCGusVdbJ5LmrOSZT9m9IX3q9jfWgXkJK
MN43R8i/ubMoFaR6+0CeFgsedDO1DnLHDN8b1z50CxngG71qeO8cj8VFvjAUvGiV
us+I4AKaD9aXs97PTi9sfp1xBi1/xLLqvWZWpRA79mR3hsGzGGgm3dpIze+OBoMQ
2ESDKemZh4xfHBea/0ZeUHlU+gY2AWsM5TdLDEEosIsgos+oh6hpDVhaJRysXRBy
NU5GY+9yDZU7hsvkJiwVzpPD00ynj8RyePZeux9ADCKfz/TFI4wlZ7Y1pHcSiKR3
dVqOADRctkOX927kOqt10eSlC4qKQ01ZhJR5+D9/Vr/nXN8UitlZoZ8+nQqydY2M
fef6r4EfDIN1M0FFeajHp+hufs/BFMiwWg2bhTAtU4i9sVxRNFmsSEi3XDylcq2F
f/LfdLxwu5R+clMBOVo7oTj9mp8a6WLmWzCkixbZhD6IfulaGG7rGAtDIXQDTSla
0iRq+15ZgkrC6jUxVn36ZNkW/K5ZM2LBtpeh8d/BViX5FD+vP88iKR54sbslguEy
L8jVie6OktKQ2nRZLF5iSIAR1gmOEDuLcVucWVRqXvvZS83OP+Z4aaZW1hnl5wce
JfqGAJz/gU/CNKVAXf64CDscmn94hf/P1jCVWDXc+wwSbJeY5NzEEMK0UJ7gbbW8
IGkVGNHwb9qNlJvWqD8tF+rUHKzg7uRSyJ3yYHIcxG4S5jNtfgxIXaWL3eIwl5NH
lUNtVceZ/qmjX9xdxeXQG+1gYCvXlPP1bS0QC+M+glsufwjeELl+lsdnoOoc7CcW
/aXwtIxKuNH8rwDBWhRe3XrXSV5tX/M/3VaS0r1UUxj4rJjm0ekSLSrIAqfol58Q
oZ06XsoODmdDxC0KdvtWTCNst4sJoZmcyNLP0w3dApyKhnzpTdR1n73CVCLfewYd
IioU/+U/FV8RCSbVIVjbn+IUPryOWirGKi4hL4ZDlmyQyFsQ1uUBC7VEJMvzPSER
OZkhyIKxQYHfs7IvynECkRf/KV19vy5FEAygaAN5VYbxyGl28mRN/JGKRo5j9wbG
4+2Fs6yYi8gnn9c+nUlRQwxv8EwgYT7PxuDPE8YPL5N5bqTV2bitgLiY1NRl2XCY
0bOeB4pYMih/SAxyz6rZwa3jaw07Y9yHzJFqc3NboUoT+oKZdnNgFLSRsfdkqGL5
kDLPiGJuHndFuEufV34bIPrcaG7xIy3sen9rTXq90awnMIPTk7Ay7sb/O1sEnACv
pOxKw7CUh6AW3sgIS1HKFhic7PHt+9+oofGWnXDGzPkAaIPg+vT9JOHJFYZY21MF
YiLuIO3bR+7Qjo+m10SMK3jtTbO8PP/LCCSONPxYieN73OYuaz5lVz4igg6uDzKr
1+1W2eYfxYModDinynp8I4IBRlMTPUBRtNi/jo3qtm8kpzvBOXjbCjMWDnjzP7Va
WMBATVLi27JC9zOMB+4qlwEGIxSC91PNy7oggiN8NXLZswyVt8J9tZ8akYIsmMLD
t/Ao3hfVKl8tSpvP0uJYF597dJdyMpzC5mw6FZlMbQxrzA3rb29sH7tf+5fTUkWG
Pi1qYKxHdPUXWhmVf/kGlXmXTXkCozD6X208omx2PQWculjjkTC0SdZtlYpNTM5r
/XWonS9p7p7/fymVkII/LebKzztFImLpLIRKp3vFdn9oDJEZfyjlg5EZlHaUr1GU
d84qxmKq/Dj18TaGFdZZBAM0hwgjaIE0BkAaySDHi6TXt2wOTqeYM1Gru6M2+ISF
W72BaKAZ4JNkXW1MpE43vEAXzhfUD72+Xq6NB5cZP+Pb814II/8zrhO2FJZPHmt4
Y5vdkEfGFB/mESHIkPbz5ZXahGJTHcUapFAoAoJPAPzPFcLvwfkvsw09EyK1uIZW
b+YVMf9cxqG23X0vZQFe6+eRXgmkKXRe7+0dGzM0BRt/5rJtCEx+QQTjONngMlWc
AMluk2i+yVDFCC4DsJ/v4fz3LwDoPQgm2SYdRFFD4TOScT9PwmDMrtZUpuyYeY87
ryuNhiwBuR/RzPHxEpn19fDHudYbc3YIjSpndO0Rrx38USMlT/YBuNim6BSw24Aq
6NQH7tUFNi0aZ4Hc8+Nhl3sxiFTyXlfh8BMop1/qLtFe2QMqgpiUTGWkEucMwVfr
L/ZgKRh2T8VK6OwTZDvphqZsVmjwVefWN16OSANI/7mAKBcwhstY+VR0K9nnzSM2
6N+M+ZX6Jg+lNvxQ08HFrb4pspAsr4vZNUEuzj7rrLbWntne0OzC8w9DGfqSG8F/
P6YcMXc5WskdDtNVGLyhCdnAmQ2JebTpFzrwv+PzxgI+o+3moiwfEo7kwyWr4OFC
mBkTJcLYuglKcygP2kB2fOcKzBFnEdgowvH+ckppy2iURHcaSlZHcqUt1z96nLU/
IGIGGDdfZP1DRYAq0PQujokcimoe4iHUStMXU4oPdJkSUz5XWaX7/66eln0C6PXw
xbOqzYyEFYP9WsKVY1n5+M46kkJ2tqft0D/EFnNqtsKbpX/lQUHP4tqVNV6SesVw
+nT8QCvznVuk6nzwbI1LQXxcnsoSf1M25CFv/2LsfbB1iMHKZvcjmGvFfSF/3Wr4
qhHp88I0IZbEjoBiYF1HYeuYW3t42RnZnXp/Z5NUodgww0qIbaPMOKAn9UqPG0dc
z5c7B1vsRhzkGMQKNkicdHPATmlROba7ZsK6oJCTt+JtVmYlvH26K/mHaS9i0zg4
+z1l0Zd8cRAPatQFpv0qL2I0CKbNMlTMUm6God8uyDbgRf+H5nlMnAlRTia0bQU0
I792y+05YcxHSzDeJhP9q2kHtsG2DUMtgHGSSL8uwF0=
`pragma protect end_protected
