// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
`pragma protect begin_protected
`pragma protect author="Altera"
`pragma protect key_keyowner="VCS"
`pragma protect key_keyname="VCS001"
`pragma protect key_method="VCS003"
`pragma protect encoding=(enctype="uuencode",bytes=200         )
`pragma protect key_block
H]J+?Y]P MRM_@3>6?<:A8:C49>*/I2P$D1>1IWWA16&H7X[?C_O#R0  
HB'UFYYI$[V7?:7R<./J8NGEQ*%I<L,$1%PY_PUQQ[T3,F7F>NR:TD0  
HMYQ=^>8B"!%N!;0C&9"KFL\7+B!IY9<RY;)3=(B\QFHQ*(*/8'SJS@  
HOC @(;%KHE6N6,29T/^#0&2)1-7W9C;&!THLIK]/T T+[7I]<WBFZ@  
H'II,#NIQ\[(@]NCT^2/)&TTX:I)8M8E7'IN<N?<+N_&7J44(;Z(%#@  
`pragma protect encoding=(enctype="uuencode",bytes=17904       )
`pragma protect data_method="aes128-cbc"
`pragma protect data_block
@D< RP?U'$=<8^0U,EKH\O 'O:P,ZT]E!@L<"+E%@,2( 
@ &8#W=_!]QZ+7<-D>KP^L. Q8_9%H8R!BME#INK=.(L 
@G++&C9)W5?)DI3)P1/:!;IB ]MO@VBW6,+E8>2 \RIT 
@>F$SC^!/:A N@Z*!I!TJ5LD]RGY4W;L12C3DDGX)2I4 
@N("WZ-\M\#+=:.XKT&O775>@1:*DEXV?Z\X"J,:680L 
@>'T@VXM4 +!] N[H*E!DPP'8R)<2=).R&6]SJ<9T9(\ 
@]8.':4HQ/2?=?!W9/&8=C/('=P:M,9.$L\68SZE+,HX 
@#WO2$+PZE+>P!N^WC?L:,JG"7WWV.2H!<QC"JK-[%1T 
@!'_L6B,TX_6Q%11!_/BKY2;22X0E<;!DN;-[#L&;8ND 
@9(@>(HQ>$KK;.;"?V0$? >26.Z0@7WK))SH*3OM+."8 
@+>M%+2+1R10K:XR>3_<-G=R.PV![PH3BWOY:Y8<M'IX 
@H%E3?'51YO*0>'L;3!Z\"DC69D3=Z5B;!@N'2HN[>7\ 
@IH=<R*]>#-_1DRO%4'AU]2--BWQF.M6XLM.1M2L."-H 
@O-&:9Y\WG:6'9UX/09":AF[QH.U=R%DY,OXU9G*K(3T 
@89)7'.H++CWX^)^?./0KFZ WE_U&.VP"G25)1WY<,XD 
@-';JC:$O:XZH@2*>J_UM&(_(P@JL6=3K^A3U"VB46;L 
@:;(50RG=-6V%",FR9JUQ,WD3'[K8^X+V2$?,0Y7ULUH 
@AZ"'L-PD72$\&B)8X&-J%/6)JJ7'6QV0#(BZ/$TL'., 
@4+<H1@5VU'4@G0LW6N5GU<XP2PX"@@T[ 4]-O7/(;\4 
@@S"TXL3_]:6,DH(Q"@T.(/7.H3P>6'+OB?).-D/KS)D 
@GS:>$FK6(0T0)9KSR/SW'X&$7J.<D=H5/JH=\*6;=H$ 
@7I5V%#H*S=M4E!E0QSA4Z6R*N*"<T]0O;L!.Z>L+1NT 
@],[N\M,3["S+3J0HDO$,H>74:VCZV-($/V>D71EB&E0 
@J2[Z<P/KY[8"/O=FR!R/.]_\=(<[MR4;-.>KSCN-[$T 
@ZVE_F X@47#DLG8ST8JK$SQN]'@D4I0.!4CT7P##ZR\ 
@>8FXI0,=[]96C5C7,N+E&/P!QKOG^OVMCOJ<\1!6Y\( 
@W9LY;9J*&UW.LPVXC<D):PPZD@VO51&YQL(C<&&.!7P 
@&OG$E:96V$;D-UEC:A,KRL [##VT=#X4Z91UQ!MEG$P 
@?-[I T5<5)5??78]@XHH+.RBU#LZ(ZN(7MG'0:3@5W$ 
@/<U5Q=J-/#4M#>.1$9S%N0K@3V]FYM6'Z)L'(;.MH@L 
@FQP9! 3$<*FE"E%VVP6^K!?9UE5ODBK4;DI%DQ#JI,0 
@PY)@%Q:$?+!PZQI,,7\@N&7;YUZ<,I+D3Q"%(U+?V_( 
@'.E4"H9D\"KGNF=O?@[?M21K<UCDR#.SZ'/R?DX];RL 
@FW@^KG3W9P1V.N< ?.=B%8(C/]#\0UC:6;/W2GBHNB, 
@E/@PP,OK=QZF/ISNA[I":Z+CD$>SIPFM(*Y6E&"A*O( 
@F$\1I@Q(^64!3Y@0//NL1:/%L=$9";$2H,>>$3P!(%0 
@^R4BD:54*<.]\[2\X[>!EEK]KV;QP(CP>;"/'/.TBC( 
@LJ- V_9$4J?6 T4>^ M^YJ5OR_/>9D)8JZ13RYBVPCP 
@$N_H4>\X*"B(+@^G;=4;+>?TRH;6F;="&?,)U'A9@RH 
@7WI39Q#V=_:O?RWSX!A,RSO 1"H.!G\Z8B@R"V"4Z?$ 
@)KG[G)4E-BI.2%!XX)Q%XV-[J(;O* 72&KKIB7D?4!T 
@43!NQLV #W/)>M6>W5^'TNG5'!2&RX.V4J*]DZJO%_H 
@-5LA=EAX]ZSSH0,O"%#J#<>#OS.#:9NSB68H&YJ06,$ 
@B!\VAC:?0HD#K;!!1HB8+)L,W&AK;U7"/*]"%R"K'(8 
@R/%%3>5A..;"4"5 IH4!JCF";H*Q'1 UK#9 >'].K(P 
@TW$"?2]-F"B;2X>V1+?(0(;B%)7MB9.L[W4A!8U+X&0 
@.*(E5JU,&I.?'QW5!##[8B3;OJ23H"PU/^LR:&#>.]8 
@E9^#1!CKR*TXL,V-8M<66X89.["9M)APB4S>)/W1PUL 
@L8W9AL"3&6U":CN8>^B-Q<BKV6$<3$EF=.<?/^R'OM\ 
@UQA6\6;/)7 $SB,I^G5LMX)3Z6^E@6X$Z:Z/!*5\S\  
@_3=9%*=:8H1^Y(K[@6F<BOKU@P=N0Y8QBG1&V(^X3(0 
@8*F^ 'P_]%WU];BN/&)WN\AG'IGJZ\  (WDA^(:&*]8 
@/IQ['4C$S6#Q[41-0P7"AW#M]7B2^S2XRGP;%2))+$\ 
@C9Z-'H[\=XZ*]R#/PK\:F*>@<R*H*!_+!&[0U[5N^:8 
@@O%EC2OOKO&B$SALGO*[V9U6>]%4O#,SP6JG)RSC6X8 
@%:Z/3TJ%DLPJAN"W]/VAXXS$,H.B$H=#@1TXFB\E0*< 
@F<P'%.YI_8"QG0@ADJ$@#MB'!B:.,)A1 P4WS8;5";L 
@KX5,X\1YWED=T_V9"*:&5!V:.Z53K.!;M7R\F!, G;@ 
@XS!AXFW<=Y:LHOP_X>.J<12RIK^#O%4M \@CVW$G0%D 
@K/)*(R[J@6V\QC>1O 78:Y\!ZD<VB(JI3=WU\%\.B*8 
@W]+SX#KM"EK*0MU4_\T"$S1NH+GD;IDWX%Q.CYP?$1L 
@=$:CG4@I"WMF]"?Q0SZU>"/^RD?RQFC=%5?]JQIW5@< 
@K0X6%KA[^06#YR(^JSX6QY>+'8XF-U"3,W]6YR^[L"P 
@1!3]41;EXY1XI^KS3&HMINK/?)\Z5U@&^+>ZK1>2Y-4 
@/]A;O\:&% T_?!':"T )QB5H7^IH^=U3M8A\TMZ&\V$ 
@@]O%?#[8[SO"Y(B9:,GX.G]X*HK=9Q\2J3'::J^9+$H 
@&V..%.]PNU'003?/Q9FRD'^D/+:EL?%A?H2*_I>$./( 
@R;Q1$?TXQ]#H*[P^X@%6H=I*+5#!V!+H+2X6Q>"6J ( 
@B#($>4EGPO"BW7(\O\MN00OMEH!!G*KT-O38D1B&ZLH 
@&6VC9>GK'HJ;=U$(<RA/@H+HFNU7QZUHQ-X.2D3*AYL 
@#TN"Z;A4K2W8:-=R+QW%O$Q@[2N"R@^@G4Y32NN*0)( 
@@W[B06@X%1"#8GF;YS93O(FMNI]54AI:W:K=^T6L:<8 
@#EXBA+*^:.2!H=P&U[L(I49R?M&;/-[=R!]5"/=NY"X 
@A)=S]$5MT9#AYW,X"G( 5D$/7'".MN@L;CHJ.X!!OQD 
@)I8%W\%=R*6D-VDF*Z(!M)/4F)!X4LS>T0NK[$DZ\*, 
@KVR'(R";)MW"BFZBCD-5#O"?P,+R^68J!48L3%E1'"D 
@PO]:-V+T44/C$,''^$9B/X54:X$&MM-^I=\/.8^U1Q< 
@"VY#*GYYBRHK!YN>_%^;!;-OCVOS7DH*(/6@5-0E:C0 
@V"_-"'3WZ'V>L%H@F-XEJ!.I#%I -]I_&S8?&T%+Q[T 
@QOAFLK?;[@A?N^B'W(0R*I/2RJ%?L\GR?V$^2ID37.L 
@R-[E^VZ$CT"&<*SA3ASPYD(_YAEO@IX!\0W(1=K@%,H 
@=WSS_\2);U<&&&MYZ&AG.C?M9=97!@/\618^(3MAT;, 
@+/^Z'6'MO*K=2OF 1%?/(2A[)I"WVB4;A_B49U8S#^P 
@YF4"#/GCF9O_BH0Q\?1<4S_ M<I&&;%1E\A>U]4BG"4 
@^]*AM66#:]6J]=FJYU]%2'5:KMNI@/FM(R!P9"R;GAD 
@C0#[)RW5.75:N S(\<ID$4&E,QD3#0J ),=&W&G/ QL 
@BHA. O-\&4:G;N:$4T;F-S="'XZ+3P<$K%YV ';W1\\ 
@#V+WWE67+G3P+6F=^%.ML7A,SZ'6F<?.G"8+"1I@KGL 
@>L%_<DU<1UM?/1-4B#]^/E*8&VGXVMTNGY7"/'4UB<8 
@)[,&M)0)X_!C19\GH/[>($F/GPT^FON&+;Q<6;6?E]T 
@51I,M$8YVGM$&%_[C 5<W30W!]DXREV+(AOS\+ZW9OH 
@MCJ6/TJMG*UB_3^WXIW<AQB2J@XO&H;XL',KY2G;U2( 
@#N6 ?=V,L[$NBPMV.,>&$ 0Y>_"DG\-4UH7)Y@@7=8H 
@<\T@J][7HTM(]%<09_M!RHQTS!'IKL9[*O0P6T'4'9< 
@D<VK+ @.'N #FW)\US!S%-]^,F>[Y>U9T@(VB.)TRWL 
@'A" ._V$%N?*#E2;MHO@I-<E)[N>"LIS-=DR7+%$8X$ 
@ ]TEV0UE5;'2RU'^AQKRZQ^KMZM]=)[TI"ZBVV%\=Y8 
@V8&RL))J3@R .I9J">1<!%;/=P?*91K["'NZ5VH\Z-8 
@?=H4L!5S:H[4:[>:4MV9\W0"-UMH+_1OJ/6D/^Z65X4 
@5I7LJ.MQ3@6#-OP!TI*5Z%G'/K'-XM7)H]Y&O:HB77@ 
@756X^9D\S,!V9T%:![PT&(?HG$G<<'/;(B/)U9Q#S)8 
@B:KU.O!*71I_2-*_E$Q>=\(*PF5=^;1+RU(73 CC7<@ 
@6F')<W!Q7"\L3E&,4*&5?"%4S>'WTM!C 5Z9ZCWZ.[H 
@.41FN+E1ZKS+8BI^!%N7)3%:Z,^'?&A+.SH]]:&&@3$ 
@HC:Y9B'<G (^MH/-[,X[_6T<3NXT]%\_@R$&"PZW1)P 
@]U<KS-2HH0B).OPK=!E+PG<D#T6HS^M3[-)!=..&(4H 
@7$XB'?(S6 #=@IXR380+9LDP1NX9O@@Y9W<GOM!:R#L 
@V*#$GD*JY:UZQSLE>Y5 9K/QII5(1KO+*^!YK\=ZY_D 
@$K(4(;E3 TD)6=D76>B\OG<:+IPB*!R'0H/DK67KBHP 
@EW[L\1=Q!))<@& ("@O"DREPP3/58=9[/77%@A$S8"D 
@U1TK4MM''9X,>+ERO!#Q6?PM&/ 4$B>F).LA1IQC@M  
@(Y+X4VWVHK>5GWR@6UJ)-X[6[V38/H2&I?G<P5[/3BL 
@OV;=4X5K$7TP[?E1+2>=LL(WD#'^>^>HR%9">/,(Z9D 
@'TK/[6X2S%G:ROC/N?/!@?]JI%3O[AV=2GM=P!NVB]< 
@M!'6S=3U?1&62JENV)D'^6JU-%W<\5#8H@-,NF$SUG$ 
@:D" 7/&.,FXY\[($6C;S26=::KVT7/4C"<@OYBXEBV4 
@B8?/W@7Y$5UM,/\2\WZG@DO/&6_8T:E?#44;^A;3W#D 
@MK01RCNQXUO)SCT+F)P>%R>7'8[R&!*&NVQS3N\HII@ 
@URV.>G]XU8,VL4"PW'/J;:YQ[6IC@TR(1EHN# @K2?H 
@39P-D;#[Y ND%GB4L!/GRYV3)M'<7:YA ]CAK'_]RP< 
@H/Z!F[+FU4FO?H5V*2F<JKO\H8(CHPF2V'.E[4+[/!P 
@SQS8_^&"V;D&'"NH?@WX_JBIR+(!&O?&D+Q7._H(,M( 
@+C/4 Y7QI8DA--]CD;4@@LG"I#IA/+?H8R6JNYC%9"( 
@#-E@?$%9>'.0!<B'Q JR::Y+:B0>KKWJMN'SX8Q(&V< 
@#XD<K?]%(Z!&R+R+0G^FB_4((3I;<]:NSK/[QHK?F6X 
@RQO63/)BQ#AX">!5HPM)9VCER7-5A@3:AS!DU9H?VL$ 
@$<#K\0OI['*<5[^)MTT"UV^9;?[#Z9Q'MJ4R@>_ZAT8 
@6F=K?<:$&%&AV/>B/DOLSA-3;+.SP*?F%U:*%E0KG(H 
@'.GBL3'YW2]?ES4(*3A%97*#1SD\.KU#(Q06-X'38KL 
@N/I690YPK;*6ZJ,!(X7\J0N7*3K*A+H!L\W8\@%1#^P 
@KL/6[EA9JS:Q=M2:4IM?86D4L@DN,UF!1%)XEOYSO#0 
@-@8]*5K4YUE=LJ5 1 W^"+"I7JR/[Y,+HR:_K&.#H:$ 
@,S1XV.TO@&"QG#0"_WP0M@H#4B<OIL#5F@B27 0 2>$ 
@N-F)'5,[2<M!S/J8! T\TZXE#!(L!_39(QT_]ND]K.$ 
@Q0*V/<07EU7;6</1PDF;H(62UEW':_AEMWFJ)5=4]9$ 
@'OS(4.ZS20X!@Z/Q()O+%QLUAA&,.9UG52(65V;R6OD 
@1*>QV#^^\5*W1".;;MOPX%%Z6T5II@ 2>;AQ\'^F# 8 
@Z&N/']_PAJZ 61D(EV$&-#_>0&'PQ?VH'E1LYUUP;*4 
@?%1EI?2JD: ]'>D@FI#;U+/Z7RBP@GB40Y+D,'2Z\7D 
@D7I).8 Y% +4BS!^:D8Z;+Q1C?_)(@=["((A@4)_BS< 
@-&U/A):9D'N+#C#8J)0CA9?3?7WD[;/H&-E6/VKEKRH 
@";. WW--3-::H^+%TP!1+Z=DI5WF#< -EUD4JRE#0>4 
@<U(EGF!CJ00/(E%M5Q/ZOGD'Z;E!$I[ZX,\1=10&L54 
@)Z9J75[5#(T0X!V8?!6._FV(QWHQM59)$Y\\*0BZ RP 
@08(0:*_')HN8.K-];)N* ^E96I3!'FX5;9N8PSSP_<T 
@1)]M- U@FC'B6G:\\!=*4+[D>:0M[J$80"A?T"W?VX, 
@0P*1VWNT\"Z$15"M8EY;DT]#"2V4VJ( Q>.A$<J^=Z$ 
@::\U>2N17''29E0+Q2*5C,$-Z+,13*NV3)ZZ&&:FT<, 
@90&-';$]Z"*A]CS%U(#].,^@M'2XX1"I;ESS#\N78C( 
@_.U$!3W6JN!"2F@K"KB"M<V,--U#D'*2R\6<JO43LW\ 
@U6K>7O'QKCR3 :3KPF+[Z%,>F.LLU 3J>UF:(^=D31X 
@RF^[/$N7]K[ZICYLB!\09EK>T@6XWZZ#:CBJAVBUX+0 
@M<]!;2V=%E:N.Y$%7Z\))G:H?"GK$@!, ;N+M3X5F4T 
@E\UJ&-Y3)&74(1S/\&25A,Z[0VW;9PRI-U._V1E]\]T 
@2/ (;++/#,:Z H%MN]126%>PN#8<6S;'3:<F%LZQ$*\ 
@;76U,&6A +;/GRXJJ0X\9R 5U9'&PX1CQN,[/4NTB4\ 
@KC'V)$0X9H;'R64XZNS':[."ZX^("<EREP==\UOAOYX 
@"I2JL^FSXV_!*JPL2^?5:J(<)5BFDEXZ/*PW(,C$)&  
@P(EJ997&#\['5)7MS0U!L,#4G]9M-53CWE!B7!E&P:  
@YMD@-C9=$!^ SE61&RY<CU'JV!RM [&N;J+$F<W27CX 
@J!%E#\9,!KI'Y4GPQ')/[H I[F_/109O[2F/+^(%+$X 
@\?43 D0->IH+8H663!$"O;N=-AJ7[#/YNR41C@(Y,[@ 
@K_U"IL7_@1.:S>JQ6OB!O@ (/"?I$),>H_#ZMC.'!'P 
@L+ S+7+Q<E]^W<@8:G36_QL!BPOQ_9;44=U?/QY:P_@ 
@)(:6V9&O,,U2B&J[R57JDZ 7SR=^<><V6*!)O-<L[F0 
@:FM$GC 7TT!PHL^J<%J*S\PM<78;U51?ZT8EARN_/YL 
@M!67I+W)6?2/IX^$X*23RJW G*CK2S#_TMI:!L(JK0\ 
@Z3%2UM<_<9"R11%[\%@!!BX+H:V("=5R+9"8QNG]99, 
@I^MZY:1PU_8#O^7IE$F /".BWC.2X<;^U$].WA$9<%H 
@(1YV  ;S;(!N%@ A@)_J3J)LBCN\N?_^; NJM>I_Y%  
@MEHX7MSBQD&I@GUY J,8!P2F;TF# +OV_NU$DTHNGF$ 
@A,F;F:B1U12GWI]A[I('"P_GAR*Y-B)@]LA,KYV=-]8 
@N6Q-[$]=A8^5Q (<R1_K#XV=UR+81^G81][J+U!9HYD 
@[ILH;Q]!WHJ$MC\S?;B:O5J@";;[>(B,_/_0+C)BCZD 
@VU B/]%O4.L%&//4RH<,2^F=81>ANWJ98U%%/:E-L'4 
@XIH"SI7?<CFS[]X"W0<H9CLL6_&.HL=?*!YR!=T5;(H 
@!5>T%Z]OX02'\4/2H=:'H1=/99(9])?J@S\1A]R!D,, 
@M'>;Y$$P50DXUJ(6MJE$S$Y6XJPVA9&TIM0@&4>C'X  
@>9(:Y<DZRPU-C12G!NOK2J:ENR2IF(:'+[:@0\=K I, 
@V(O6:3(>PGS[MEEF?K69[V1>Q28>^N?9'W7HX^ 390$ 
@DG/6:9%C-F/M N[,166.Q"B(CC; 'O5VQ9V]2X;%$0\ 
@46-3,!90'"<+BE)TW&M("-ETN^JSG%&@-[T0OH2?[;P 
@L;&A4-=C"&>Y_@%+\M4G>1PPW74[E$0\BN@ 4:+DIU( 
@3SY]S.V)E2Q;# 4C7[[?UQ7>67;02KN,<#'$$E#6D7( 
@;=3;1IH0(#1^%+;+WT(^V^!F=36Y#1\J4!\**#F1RT, 
@(L8;(V]?(N2GL"^PXK@UO$1T&75=K\=[^NK7\FWM/1( 
@&E;(.R5 HZJ-E#]%O J#8CDQ^&22/*E@MU](EY-U#24 
@_H)Z#@[,6-<C%[/ 65(KFV>7<'Q:RWDQ.VFZUYXRHB\ 
@RU6(C$>N;LR*#EJQ-XOEK!#K9XXF&;9E^3B)<ZBR@3L 
@(]E@++'P2HMT"8=J+BHZR01%=Q7"I;)\M4D[CQ9O ^4 
@5T%Q0#"I8![A%36RC!:$8W&_T0YQG=D#J)M9]@:.92T 
@<U*;CM:DFI?#TIO>=?SH<0AUI^L9V_0,WJ+NH+6J74\ 
@R?T!4R\RZ&4%U:L'5>1> 9HB;"SS1(QTZ'PY7)S=3ZH 
@GGCN468A.)<?HA:$T?Z'ZFHD.#!VO'' P9+Y28!F*%D 
@:I\4O-M/54COEWL8B-/_@';=>Q>0XXD4U#4#*S71B8X 
@62<7ZKBB:.*C(I$7%]^F.MIA-QH!,E,[RH2/9.6:H\8 
@@/LW=8$MYZ%3[$9W=9W,<:M-"QR@0S^H.:^[Q9IW+!P 
@ K28>3P2723\]##@]>&15]L'M5T]*G6_X6F B<P=L$T 
@H*WTDZ<9:@VC\X<%-A2>NK7'5F:,%+3T'+U\])WR,F4 
@4+?IEB#^**](J6-:?>@GXDSLB<F13PK@!FZZ@1?P4]P 
@/OH/AH3HNT]$DOK)3_O5N$] &W&SM4'7^SS98[7:P>P 
@^ZQ0-T+BI_[[A/+J.& 8%^O#EX=W=B#JE3,=@X@&258 
@F2'PZ4<%U62_;H>?22^+K<6UFJ##PSE$=1V,/3T>1F\ 
@E10C1R>,B\[D&5V\JQTJR0/"11J1:Q=?(9,/\R_XS#0 
@S&J$;1(G-KE\J[>4>BYU@']TBWT9F_321L^HA,%K;I, 
@LVCZ"$*1:>Q&S"&4[%67Z%&,U!O* ACUY\XJ16?'B24 
@A&U5[@[VK/-=!L^NY9I3-R*HXGWV2R-KSUT"7L.*@6D 
@\N]VKNGZIEJ62%W!A&&]@#\\_]@/@UQ8AMLBP(C->&  
@W=L:-4&Q%;8]'&0&>?$!K+I25&&/QD9APMM41=,HV.0 
@'9C[#^6]B8PY _^W_# OI'4[VL6$@0\G<?T":-!]_UH 
@K)-N+$=<%'-B%OR+C6L::JW5FXD2J%8_(K1Q*X4:3K@ 
@/>MV:#:E??+D3B55J0*ZK=X7OB;1A6,<./6"I[2P.UT 
@@UN<Z8O6$^L00#%03?IDJ:"'NA[Q_@\\&'D)^"JEFXL 
@E(?D?J%^GLX#;0%!(7!_4Y?V1H+;"@/?MIHC[S(U6L  
@O.OL""BGFA,C<P]&@U_!#]*4()TL5-([D5?%O1/T07D 
@&P&M\687-P6-FWB^#M7F4@^Z)U?)/Z#0.7S?J!M VW0 
@)BEH>I4N@D5*T37YU,5!;;;*KOGF5-X DEO8ADE(B<0 
@?X<#-6A[7!I#'7XA-S,LC-:_0-\$7*O0E32OXD5L_<  
@(P%7.Y$MSSS48N]/E_+Y/IW,YKO.OYWX-M$RK^C.6F( 
@L'^/@,"087^@7Q9_N&N&@IJ*]Y?=5>EB:243VF ?G?@ 
@4L7,KIH-,O\GX,)4E-GQ#-A]Z?E8EZ>G6Y91D1IA$D4 
@>,*R>JFMT"^6$"AA(LIC1<EX.Z?ZFX$>Y?9?PR==NVT 
@?Y;KU'E!,)1M$.)K1QA^)[\Q<I557P2G8[W:>?JP"/\ 
@IAN\0Q02-0-B;-A7IA1J3';+ZF7#Y%)5JE+&K7+FP!\ 
@CN .R!]!W0HK"+F,-,YJ.AM^APXO ^B3 >M&MZ$M%<P 
@Z^G+>CKXC>CEHF;(4[$R03EPV]C""7C,!V#/V<B$?4P 
@Z>DIKW9YHRVKLU ,Z3%!=X 197GS]SF+R.PC&C>HZKL 
@Z[/6DO*S+9PIGF'12A@D*)1UXB@6<BM%YE$O$P0U^)T 
@*F]2C E:_?6OE><3\N1K=R0NV!)61QVIOYC:*T619UL 
@V:14S:6$CAU07>$$366;\=JY^#W@=RH/"_3N>-_.6#\ 
@(1I\ATT4A)+T-C%AKYE520[9HO4>+C6,CYI"\-6D%=( 
@ N]*6:(N@/.Y'L]VKN:.,U2<Q&%'[+^H2B$XZ^5\R8$ 
@:13?U FS=UGA*]4I2[A$WCM\0E"F56TB?$86-[$N3[T 
@(VC077<1H^AN+=?(W#1@3]P[=BD1;FL#3.#!5L<B3#$ 
@D,B$YA!Y32'!" GC4%V"@4B#?/:Z[4L/&'L>\6]K1J\ 
@E'W;^6X \^%3GGT8L>3KM(X>HW**6].732$J3#O?1?H 
@>1+V]!.3L3U%_4&^HXG4F+:I?X=:P 28D/X!/I;A_G0 
@AR!2B+JH$ZKL(2K?HU>D#(21#T/"YR7J$]2#5. /L=X 
@78U_SZ_PQMMVPO?^>?(95_%O\I8+'B&GX^U8_/"$G/( 
@9GQ)Y[0.:/@M#I;.SN-M:6F":$7H64^>N\N_#DL@Q3< 
@97RYZN*KO,^/,L([>4%[O39E+-Z81^7QT)40HZ8:2O$ 
@0;Y;PY$8S4D*C)BQAHDH]KB2"7QF@,9AN %J9K%THZ  
@;;-8 ?3ET=9#,*Z")<CHK$#L48=J>8T>!\H4'1<@86T 
@#G;5(&DX@Z$+J&X_OZ]6MV-ZWWD&M.V0.NRH!-"<-/\ 
@XMA VT[@CF9S$[WY!^/5,A$8#K17* ^GPET4P]!=%&, 
@+I3*(I2;5=X:G4$<FGK6E+KPU5@BQ^5%=3LM,1H#8'\ 
@L,TYUPZZO0\EF_7(8ZV@9;^J^^K0C3KS=V?%Y%'<Y5P 
@4GB4+ +M]IBQU+,I4'YB7+6Q( TGD%[2VF3WN:P2\/< 
@^DZK[1V>1,_DY L'(_#C<CO(\W=UG04](F+>L]!Y,1X 
@GWLD#1ABD_&H8XYC+80F0ALY,F;?_30!/97)]9"]?@0 
@8Y$);UV,:WHLCAI=Y01AD9W%?%TI1415,L*%/TFNJOP 
@:C"Y#\XM&_X$SBP><;4#)4T5BL:G1"?"#Y*0/=#-3\( 
@9-CW^M7\=?:_(IR K>'4.@ <-*F;Y&1PT5+QR8'1N2$ 
@9FWX*3=^-C?8=(2VCN,WU4?6!Z@');DE+(ME^.D V7, 
@:EKNO(.1[ N]=^DG/X/QVSEM+?8RQY#Z[V\T/78K(_X 
@*&M _#M!4\>7?W:QT?QU-)'\X3@2_OU(DQP"!8(;Q.@ 
@6KQ7$&YD0==I<#)\[Z:VT3P;,#-E]512?_,8]"48/3$ 
@W"Y9BWUI/<8Z_7.+1EXEBSTKHG4![6>&*5P@.E:5M:L 
@3M"^2#61>]'5 B^-RVHZCD%<Y8=,>SOI0"1_G.H-GRP 
@.R>!SQMD'\(CN(R^"*NG12+P'&]:Q]V;_0"\8.>LUYP 
@59H!157^R!N%!6/8A-%O^'=XQM;!>4UKFYHFQ@\9LW8 
@:-W>_)#?R((:)TLE@>LXL'$?&*]+#_6.J[P+4+I'WBP 
@78L#O"0;:7YH,L<D9S' WS00M(G!>858*''Z$X^39*$ 
@Z#>L^L@$"]266@/XKVY8102+,L_0F''/ W'+V0P$'04 
@R8N)'V($/>0$IUM,[<LZ'.URV\D]6NE[NF1I$JD#+@L 
@<)N4\Z#$/:I0(<VXX"/G[\%&E%*[O31 M/<;72^WC60 
@MA^(MP @70:>+T(^Q?0J?@S7=JR]FW]1)\'[\C"(@-@ 
@K33_N[OR-O7U=F313;#@K:Q=%9A<<.2.F8&2I:.1PYX 
@M\<F^9RMDW-R[H&@_4<1@B$<*4,#56\W=2+ZX@8V9!, 
@V7MIU@,J%^WA^>_K>'8^SG?S'R-[LJ89IOO=]>&@9G  
@];E;A\+I;D7F,L$ 2HQ$1";>L@1'\QO]1^UW]:7-8UD 
@;63PPEA'H;1X5$A8NX JJ$Y_"N[R.D"EF$[5L0?>ISH 
@O+M!'@D_0VRZY2U3I--)M3E]B+.N*,)-W8I#^*@\E#< 
@;6R.SN-"^-G2V'AMP+X+ZZ9%X"<M<G<O?5-!1*/_3\T 
@$S3 #Y62^[NG;CAUC,D)4Y<9B+\N2/-@K +G==@_\W0 
@)#K.,A%>+QI&9Z'_HM68I<^FSW]()#H7)<]B$Y("<.0 
@T(H:)8HP46)^L?Y<D@=?/323BCY+6./3S4"F\:'A/Z8 
@QD1;FSN_=+_+G,(5=T-<D"?>I%/#8<N7S(V>X53+N!( 
@82^;R< ,R$R+I#?:448*!88%O,>BB7&AOH)TGB;WF6  
@<,3JK%*[=;>H4S=_7FJ%8:W)UJE*#=\/WHJ&](.(^Z@ 
@Y0VK USO;=Y*][/B1&MK3E&,/.B<J=Q6,^FLP!6?+E, 
@QM12^+ \1#O]3ZGZ1&$N6Y!6H9+7'%_P08/9;XO26J\ 
@E4"N1CJT"IQ;_C<[M6:,^Z=J'O]PM!4A_+>YBC0)1&  
@"E?YH^;V$JOEHI'V6C](/2M'>6= %6M[TA(RP5\!(7H 
@1=S-JKG^?GL@-Y?:#%BO42.UCY4T)C*XO1I3<OM6:)  
@/@L)6>:E+B]JP[O-YSU(2EWE.J8%LJ!PIW5@?Z$' /\ 
@K&,U+V0W<C[Z,B;Q^L^KR=S;'DX/#FYP)UEM &]C03\ 
@M++K\J8= V!]<Z&8PO*1J.>?'J2OX5N6))SACYI17NP 
@TB24"8/?R?#[&RMY#\4)L\^]-]P +L9E2D2 (1NQ+>L 
@V_/7$4/O$ T,E-[J/[H9)/B"$ #GW!,K33T2+H<DF 4 
@'G;&A>.4@7?$:Z\ T5LM"8&NW(I:UU4B%>V>6,5=ZT$ 
@)&6WW'W5^@D85>7@P3F2U,XP'KO$J_C#?B]QB$J@NX( 
@KRYR X]&_>PSZ9.+ /^=;JU?9[B=;>G,U*XBH.R56<P 
@H+P5BE*68]GB';FR]SW<87I/43*QQNOD9$&U\=E/.[< 
@6*HL9 :>01J?I11BPYLQD"NHV%SU$ T1R06N&H9K)>X 
@Z_? )$014#6W%Q[HT(W=P<H"Z$Y9 ]KUZ+WE1/F^_Q, 
@%@GM7D\7Z0M>FUDWY_V%\UFX@WF3D1O19Y6YO^;*BI< 
@\1$I&FP9F1S()W,>3'HU.P&8B&N$"#H4LC%!(HK?<+D 
@_9YD\BJN57#:#6HFH=W4JNF;DJ:8G?+R_4SZX6K\B:  
@H3X\ZL42I [LD7+_9U(@%>C6[)R_$#.9HLN;)Y233MT 
@*L\%V/4^\RL6R-]ID9!!Q[WGOY)#E03*+!.?]:([418 
@[T'=ZSRWS\<^GS[0H.8?,U]BIZ>XGH8%9)Q:(;Q[TP@ 
@:;U<*)9\P[88S3*?-(%K/M5K(V!Q8+<(I"@'N&K>F!H 
@_2!^N>3+,$#LV+R6UAR'&\Y](E\ AJ\ID4C!??9_=;L 
@093Y,IN766P?>&5.B'&UQLT[P_DBYZ6I\*B$@\)+$GP 
@>!.G:TM',U##!V!Z[W#K3Q]6(,X<N+<3?$^(*\YTQ-0 
@9Y7^\<.Z4ZD&$YGI9R0<[I:GL=3T@2ZUZM@M>UM:^A$ 
@[2ZT1!J7@)"F3XV2<W-ML]_20BDA(HX8#TZT*+O@-+, 
@H3LQ[H<[G/8LDV.&Z/6A.0,91#')7DN&]=#$:('_,3, 
@5\B6L?<YS,-O.R*:212"WO*CNS3M =3@['%O8+'7HSD 
@.2GMN6N!X!R@N,95-,3C<4'"N;5Y+ ("-1]4+#%3D_$ 
@^AP)$9*!NR*(\;,TNLZU<U;[:HI:D <VNSF^IS8?BGP 
@9?*HB6O2Q,LEGM$O0$5WV1 J@<KMHG82N)XPY\A5[9L 
@79^RP1:78L'AK :;&LHW'=$P?8GW>M2SWC5>+"FH)&$ 
@X$N2F^/I?+<+7OCNHTOW$.4^Y"9.P:W-=@Q:1744A=( 
@8&WE:L/\=K (>-FKRN"- *=R28QR"A#+M\N2US9"^^H 
@,>GJHAQ(GBPL9<C^W4<315>5J>>/G(UT=>PD2$@H-T$ 
@MW1G%GM<0)T+__P8N+XF$X(&(X-@EM:X7CM7Z56-]=\ 
@^NG]".NM#+*(']+<%GE])<?L%[E),0#HL*>>O6W+L90 
@K'=,,XF*L9PII9L^%KYO4G-FXI8VS.)+C R>@)QE%4X 
@,V7S;D*HD'N:B/1(L5CY#9';YX)L1,&/2(EU,".1?P4 
@5A5?X.WVK7@AIP45E2^5QP2^3U'JXF\Q]=" 9ZD1*<( 
@W/?/D()?K3K.):YPE[6+' I<,BXN$MFN</9!P>SAS1$ 
@2,4#0U)5J,J78=Q:8?W!A1]D[CIC>U?OI^W:[&F-_Q8 
@O+=S'R]?2L+1:':M]^:AG9O/9W8$%=G4'G'5IQI,F&P 
@S2$JQS$V_,;BU2M ",6#X.98\%]4"$9AJ0 9=KA8P6< 
@4N$-1,_=M*G@GZ[F0DB*[DB%G>NM'AA);X:6P?( ^$X 
@/U(,@H\O1,>-?U='3@P$ DC5!^OW_O(1B76:.+/$2VH 
@* Z4<ZY&0E-R22:S\(##T'==!=*.@-E<IBE]]P-7H#< 
@VJQTE+&'A*5210#\BJD<;X;X%(3#L%HJ_=;#+=?ZM.@ 
@<=H26HBPJ4L6X:"L5J!@].%FTT23&VQT=!Y;;/].J)H 
@UXR9XPLM7##)C=RG-4&C96:&H;X=_#$?2FT7F6!,D P 
@$K"C;#Z3*$/GN7_U"1\PR!:"LSF:@;FLV;?-=P64PW$ 
@"GK)J04SU(6@Z.WM9B;FC<^R3;EH2V]!^BQV6@> <F< 
@(Q?^(XS""=NL4U0JR@UCPB@K,&>4_-](K<T]6B,"<)H 
@[ QT-3KG<&K)15Q+)WPZAV+!M%[]V4*]J_N%SG5A)]L 
@?TEZK.EF4_&<W.>.EH2:3.D[U-/XHE8N7F_1JY6C^F4 
@+XQQ4:;>7A@24B1QB[>:O6M.,]=S"-@C [C*Q'1_+D( 
@C4-2(5[*59Z7(2(V["??4!A1GW"GA63:_ZE&]Y_C/[D 
@6<[>_P>%L&>A_3Z-ZPRTCL94SK$WU;V+0'O7#V)$T3P 
@OR>X5P>VZ*<Y6]PZFD.:>5_W$A+= 8;209V/9V#Y&C  
@UKIKA0,FV[)MHQD*#%TZ9CSL5_':W1]OA%"3ZK6ZF#@ 
@"Q'I<<VO4D;U#.:B8Z GH3"?20[)Y:C?H.J?C^GR(_H 
@'PBUW.(^I&U(VD6=.H>,9G9Q+UI+.0+!MYNBE=:U5\T 
@Z)TG*5X(85W.3/S&2QU"_BH[AFU%J%Z1!Q<<4*]6!ZX 
@M./\3;>D3-CUF4P>LR$WB=\V<M_4 VV(O-4#)6=*#N8 
@_CAAI_>C&I[6"B=FOU,LM9]Z1R7HE<C CFM!61DLQ_D 
@J97QI%ZA2/H>VWH82HNMU%V5J-&!2PZZ!+RY?&Y:\ZT 
@C>"SA8MX4(_&#3(.BU^2CHJD)W2WI#/9*:KFM#+:G)( 
@\!,R%UX)Y3*9R3]ORL5NJ40?9J+ <JVJB 8!);$J22$ 
@;F_"+ C(3E;_'60M Q<O3)12H54WL9MI/NU$6&TF;+0 
@S\\</S0)$STG:ZJ!<?&%@87_X#_V7\C%S%T-7;/%TH( 
@UOS2(1 $QY.NW]G93)3+ABB#LO:!?/*)X4]:9GO<YZ@ 
@8 [S; 8$&RR7E_Z"_&U@7&"<*#O;2N8O;->N 4_8.NT 
@F"OWM!W2QT3J5X3L0&DT8F$ZB68@[JXR\2-@XL_8#K0 
@B%DZ YQ= 3FZ2!UFO]Z$!#&2D:JM[Y6@XK(EKBFQ]BL 
@Z?Z), ?/2D*,_)W))/_Z/.  <[4TYJRQE<_SVV97&_0 
@MV_?\@59!G-Z0DAPM*WZE&B@1KDO2B4:,0$%VHS*?-  
@VL$Q$V:O3AC/[T#U\ZB$UW,-BD";34LTHHFZ%+A/]+( 
@;AJ/ R'60J"_%C$F(TLU>QOPS']!A]6U2LO/8FL$+^0 
@E*(I5+$ +E(LJ7&A0 "52#FHLKHC10_-/.C  ?G+,AH 
@'H?=#CBQ@E[Y,L%*U@6T+]^9 _9\B/JFP0#$CRC)".$ 
@QYA7SGCE<73?LZG%GLD;!9F9EDMR D-4G_0K:2D:9C  
@[R:.(QA$Y/XZ7[)4LN%Q$35%H!CGI.YJH0:6!4)$YJ$ 
@["T$S,>%LJZV#8!8-3&)P,P);%"<.#R_DCUILI(08A$ 
@S* SVAF1"012UA_2QJCOPM/H3+7I&*&6Q!F5VSXD,1L 
@)&9;@? *?/6IAEFO;]!0KGZ"CX:)CX2QU1;?\[ATEJ, 
@67D^B6@^E>O'@:E2 J=&YQFF36.?6FDIM#NGF54RD3, 
@,F57=X!GXC!3VC 17P;EJ57ZLTP6FG3--0&/$>9X"&@ 
@2%^(U+49:)S>/!RD!+3XZJ$RI@4WTD$8=DW0KV3L:F8 
@],:]Y.*%0)65GD]7OSVJ=G>IP\?,*B?H/^RL.72ZZ7X 
@KO$<3O5."W[<D>4BF_5;/*K2!J54\FT"OX=I$.G(@>\ 
@=@9LS6QWM*G+-1%9%W^\)80_9+>SOWLGA;KK?2AO>"H 
@E<CZ:1^+SQI3?N1VL2]#36NF!7#8P?WLV?<Z\VB3FN$ 
@28_;9@\_A90FSA68<U$S46A5E/#JTLVY2V+RR[X]Q5\ 
@MB-[*U,!""%"BWJZR P1Z2<E'9&DP\C<'Y(*8:KLG-$ 
@.0;)7D<\IV.:&/V5IX8?;SFHA][4H1_2J['CQC>LO+0 
@ , B.'6@Z]A/8=1ILH@\#5!A%DR$\(K>V??O^A90I?4 
@72D\E;RN).RZ_/*>>YPS.,ATN]4E*"3[-VYGB,ETDML 
@'QU8$UVZA_=QWG(6A&+CB72'A_@L(9Q J\J6EV@&A^, 
@\Q1<C(1ERM>3K:%:.%:6V941F#P[_-_3C#>[7> 'I9\ 
@P+ L_^LG #R(1O%NR\SFH7"/G,8(4-186:G.%/_Q2.P 
@D=*^>''_UD2J=YNF@ )+MGW@ECH%PS5B7XQ$4_E4 O< 
@03H)96L*R%,4('3!],+R[I?_J(TWIJF#WY'01='@G+X 
@N7$-8QD00(VC :IHGYR%N1RC]:</NYY/&X(("5&;3&( 
@!U!'(E1B0L'R3N,*5:$QJMG;XB@-9\$SF-GM\#.9 VL 
@HKA?%C0=*8^MXWK#&?RLX/&ZI]+1;X&;N@!]CO0X7.( 
@1HYE9"]RWT+KLI^6!-F\G0U]]II^CO]K1?CK)\B!E0L 
@\GI.,*\*!GU:Z]LK4_<E,"3T+]<K5':AWZ\11/3YI@T 
@GYI[S5*=V//<^B;#&SZKSWX81QZ\<G1W?87D.][K$L0 
@<I]0"],=W-$+M,#2^RJF.G%:R#(E3?X, >-/G*?Y9^, 
@N*9M^?U0%<"Z<*.0MXW;'[\/[KHE+5M:$C5&B*:9.AH 
@\M3GR=+W6M&,N,1KQW>*RKHTK*Q;,?9"^5W,.#]ZS1@ 
@SR /%G,Z]4C._DJ,&(Y64V.6T%7=H)B99  Y)_7,KB\ 
@;\C[\A$@ANJXD_6A\''/R:Y.?6T.).:>??DIQ5>I'&P 
@8#@-NQ_^>LYCQA  \;7@J([ ?AC@7=NQ@&*![0+]?/0 
@P;MY5^BP;KQTCVK:;&OTZS4_;>?1D@$_E >$NC^:KW$ 
@R.QAK<?4H#YL(Q@U%!A="^E_ ,:+YZ9#20S]JG?*8JP 
@*!2'[2 6"1?([HA-4HJJ4L^%PQ[:/$QXF6;8>L4IO+, 
@8/D?>H((#P,#"^\!K&:SSITRW3'-,4K7=4?<(Z+ XV  
@Z+["0H0'8_^&C'X8QQK]%+&F51)MUCU;GTV;V2G?EX, 
@X/O*BV.P6$I0VUW/&-.Q05Q\C)D&*";>!E)1X;E?J<$ 
@$[$"^LQW<>-6RWH4XH' O4-.5<,$5_L<)XJ@_!RK)DH 
@3ABCD>D*P?K'[!?S6URC-#5X L"QJ*(IK$?WLXUY8_T 
@.LM:#PR-JM0U01<<ZZ;2#<9!D*0]4 &1RTJJ(%BO:T  
@DV#G#A+KD"U:[:8A_8A(&+]2CSVTMGN.F/I*T!".C.0 
@1"? ("LWOMM]S<6'QT;,G1/=F2B5W$3JIY9ON)E,P\( 
@);Y#J9G!Q+3_][&BVH#[ZD11ZCX2,BUPQY/(<J6X/B, 
@$J6L:**GLEF^^^;[H:D4>7;R#6Q>56OR/G!/81=O6^< 
@,%"7KF5#NB,M$'36N%A!_.\8T^E<6#[S&)G*W'WX'ET 
@XD$PI9),3%'@)R49(MF(H54:UZ SRI5;L-Z)^V/?7%X 
@EO@?DC9E3KH;1U7"'UXY8DBC87OJT.=S25[:=!8'T@4 
@JL21C4<SX),F&9Z1.I,[TN%+&RSZC#KP"7!EPD>AC8H 
@"B_&%<KC'!*%? UO:R.XH.4?JT"%0"QI 0K$P(*B]%4 
@J^Y1&^;0S^_[ZIH!X02Y3@";9W,*UTI%592)QK.B0.D 
@8RF?<KJJKQ92P#7>!P,?41:YK=/$M.0,T.<.90FK"VT 
@3^QYXV?HLU5O2=[QMUHY(B<69.MM4%*>K C/JCL37W\ 
@C!DX8<*@,7YG:78<N@7\.[+5Y0FZDN%?&[^4O NL$"  
@E_8(G(;3(%Z1MX^D(3>NI!])Q58,PBBGNS'?8#>5DR< 
@ID\BP,(9P[97)0:B9 N %Z:FKT_H<6.^W0<RU'$JG3T 
@J?!;RT3*JNLU^B)'FC#OF"57>29XL3G1^;G4Y1>UVA@ 
@^/W#$RPP\8X>>^%)2E@UGL]LMXXJI49%J8;.9P6N*\T 
@F?,%7^T$FVRA?ES$^<\JH<?;98PKNKA&48G2,C52;#@ 
@-=KZ3F"47TC;PQ-VX#)$=TU^M0U"*S'P1 0CRU(QL<$ 
@- <?AS.PB \(AOWC,E_>[MM40P@D<M\1EQX(![915[  
@4F,L;H+JZ\SP34]M1VHZ&0.!U(QQQ_-;AU\=S\2F:80 
@2\Y5:*!)(7K'F@I8,):S&37-25L]-XK<;"3TB^(17ZT 
@;CORK!1"JM[;7+I[WYT564\]I;J]QE#(%XEJ,38^1T( 
@D5Q[C5B:M&;3J,VDJ'DNP<KW]@D0I\ZS!@YNX-"6QP< 
@W$VIU1+<(3/.)-0DK9WN[3VB%;1[ \] #NU"^3,I<B  
@5ZK'?")2>R;D=3D 01+P/.2G6Z&;DUXRY#- *>/RS$$ 
@19KY)KL]M%2"MU(_AX<?=="U^GO"T;CU0-U[Y7+K\)@ 
@9@RF.+:BBN2;+T#%8U6-^GDID$)K[ UM#/9+TN"S)O  
@FF]T379HN7FV(I,><$WLCP/*'1!OFVI5'OWU%N_$-6< 
@:Z]W9=:)Y JBT$/*=JB.!J>$_N-AS\2?HO ZR.50#]H 
@/4NE:0+6LOM0"87E,D'CYRN.,_]%V(RW?%7BXWCL(P$ 
@F$JH9S<^=A[+&GO*F%=3EV<1WFPP?#'EF#O:(&O&_M$ 
@]4P]95KJO;,B1I/1W7 X*Q)VEED=Y5U%@@C</O]US+L 
@7$8,E*![U/QL>EC)$N1J80I_=<B9$NBN[L8!0VMHM7$ 
@G<!JP1BUZFK.JR&)T3;H.%Z7^J-A_;OGZ.'R!P]2?Z0 
@[5=BE9J#*22XW@QH%]5L+-HG)N)<T;0:JA.ENW73\4@ 
@=$5Y_B =?6Q&44H2SE2,CTPHLP(?=A'T9_:0O0%>'2\ 
@W>!7>B?3-8!WE)A]I5+G\\P@O0=-DVEZ^4%'U);WQ], 
@Z^'9Q^-[^Z&!($Q2WL!(V^T0&_U5T*B.EUY6&0^^P2$ 
@^)'_+E<()$P-R!%YPX!!;(]-#_,0#FB>:82#IHO>J3< 
@/A]);FJVX;M4EFF#9V+#HGV7\@NB)PESF+S5?2=0T1H 
@N.N?-6<Z'0I;SO2MA$,'[)SLHZURI\]%N_CJ[D/<-58 
@,766??=(D0_]0$NA-C]/S'C?GG&EZ&(%H:$L(8QBS"L 
@2V%VC 4.@5J9/ >:?.YY%E19@/.%_IOXGRY>?)\">2, 
@%O0WU42RI3#NL-N&SA3\;&I7P4'Y&4J&,4$/WXY]R$@ 
@-1.@8XY!J$UO%67CM\'J#"4\634:)<S%O5'9R? 5ER$ 
@2JQA!)$[SX4(*"J4@[22=3SD,CGCI\F-X>E.]8$":[\ 
@A2J*Z;?3G+O;'B<?DP)VR12Z)=0$91Z@G&I&_1H;$:P 
@@.LI,<&J3A+0P_*QKZD1LBMBE]C<ID/;:_K%0T-\D-( 
@;"[#^$SK_]XM(^L"XH06R"CM>YO0%%(<ZI*L'JG?.A@ 
@K##C2Q)T+5+Z;M?ZRHY!,NQR$!TN&FB)0=,-:AHBXQ< 
@+P\/2&KNL#\<-.T2QMM+XULWA&L55GE/4XV? 'E?N;8 
@J5!(EGKT#0Q6?ZGJ4/$C!#=[4I>X2 @+JY+_S])3<&4 
@OS>A;_&MW]I)I#X?$EKWQK20ZL,(5\FCZIN/)P0NV'T 
@E[0;K))1_6T0:YZ70W3R1,,9U0'\=15(X:7H>5AS47X 
@HX:%$(;NME40SEN7.6ZR]?]H72CYUZ'OV+U%O-N;GGD 
@AWV=.H;)S^<2(0J&P0#-:.KR^()2?FTD<7K@R]_%5\( 
@ATW--6$JJTA<#%KXP@1C3/%ZVDBLRD/8PX.#97#KO30 
@B,=7'>-&(:5#+X80!9DQ4_E'5XKL L,>_@LA1_N;#YT 
@N04VFW@?J!GMK/S+99S4\.EA<I)TOG%?>=&Q@S+<T@4 
@R4(^?@Q_8 P$?S/0'\E@@/06F,HQVH0ZF(&V%0%\_=  
@L<^!1&&:4JP<ON!R:IC9S.)F2KOL^H8^F&)^E2_(P(T 
@YG9$<243#>1\=L/F>O([ZRYAOV0;<*V3FNY+KV&!VR4 
@D\K@IM>M(W5[C3U%[+MAXY$S.I0 O>V$>!C-EPZ/(OX 
@B7I<L+SO;7M4T =H_C&(L/7_EE!=>O2RK_Z48WE_W*X 
@K[F[9?$%1NZW=@S("*>\]4Z=(%,]W-8\GV0]/5^<=*L 
@ZRJ=7W2/R@;N1R(- I,B%R=KW6>L"2H/SC&\JX./--$ 
@Y,^#%2"=/.PP6ESI%Y["8#9^3>3-WPD;CM"(GB>9=O( 
@[<-9=SK^8TFO2ZZBM);,$L[+S0;J_N*]*8*[1^U,M24 
@$Y.\&Y2D=:;@S"8D-E45'%^BV.K#@:!2)I!X#*-V40< 
@G:+J$<<=1&XQ_'M^XFPW!%_'N'F>AF0MY^S5FC!N,+D 
@5=!=>U:Z0$0\&.^9,4/D=PAJ?R7A2=Y2Q(9=96Y:!3X 
@M K/!YAIM JZAB"TR_'OXR E\K_F="0?(&,3=$$A\,4 
@Q_V9R(@^NZU$W J'KR,0^VG)..6Y[!&90WE8AC]+S0\ 
@2XD9@VVA%2)%&Z#X';WJ4W2Q3M!G_8)O]OY@+:)^VYT 
@)\@&R &AKS!0]-(\E(W&;PX)W5\&+"Q5>U C:>-_.YD 
@A@^E"NH86>-2_5H%&KNW[)-ZQH5KZ3 ?_*J8%A'*R3P 
@7_?0Y>&0?B<)2*(Z]^,BI< ]_N8%XE=?7)XB]N 5)B0 
@;$K$U:E@(44Q@#.NZ]QT#1,Z6>9%C 4MK 5FY%4/ZJX 
@X 2K-JIYB[ R#"JV=MV\>0'U-Z('BZ5M6U6T#STQN;8 
@ALOW<A@FE?OHQ<@%VYE&^7 OT[A$\FTFR#/^+7K\*1@ 
@[&<SY3?.M6<'2$N?0E"UE^ST\?;E@M=\8+?-5 J1OS0 
@QW*=RJ3<2 TXHI4UN:PG 8U_FT,5R6Y"G3-R<JRT0T  
@>8P%N\+$ZJ^24E3]?XQ+<YP31H$L^PU_R@JI:\LY,\$ 
@%KVAZ\"U_T@<ZE(2^Y!XF C&.T\>+LE?S=4&XRH@2"P 
@"7K0[A-W>XJJRZIX@WF_-9M:.LVDZ//50VK=(*M0YO$ 
@[3WV%>[:JORR0[B5G!IP&;E.-P_-8KI?^F7>1BV4S+T 
@VPP5?Y>'N5]5T<+&1W7@A:KS\R\%?V4HW"S<%$COL?L 
@,!?MN[>DU:0;E;:$M_G)7D.?KXMDXS9'F;\*M^>BXU0 
@E)S';0#?-K$<\+(FVVN&2C+1NV5T7GC4^_S]L+<]O[4 
@WC/\(@OV=LQK896%#4HB2P1WRLOW0Z0: B6/#AF\_JX 
@\Z6JD=1!JB!+_U(,2=JFK@Q:?*^<O_FM2+!&:7E,0-, 
@F+FX:P6!#1DM]_[A"O?(I,[68L!^QR(:(;AE@ 4.=$P 
@I11A&MB0,$L)TZ5/,F3(TMY__)/6+%_6LU!-8:>YCKP 
@FJ.NZF[*DUL"G)J,J=+1C2Y6P'D\KIW-[0?8@E- ^U  
@KMS$GCO,4W)SVS&?/(\F__J#F<1F3A!BWFWN'>XM9B( 
@\E".P<JAI8?DZV_\A:R\#&[&,KN<0]' (M%65M)9<UX 
@>*79 <V3*+5_)WWRW^:)9YWVTL'GR)G=(VE?HOETJ*H 
@PND[<SE;(SEI(CV#3&HBP-UN)XEXQ#Y(. ?R32QK)_8 
@ <*F<C31A+#N02WL25JF\$TA+1-O;&IL9_<@1N8R3=L 
@-"LK48M9PV:8TG+NW+$<G:Z7V:A),+N@$T+_<U@ZK2X 
@!R.QK] 6D==>32ZMQ_EW!.?>C<-*/@WO-L!DW+[Q';0 
@C(:TB''-VT6\U+$F,KSQ=BCU _\IA>"-#].W*NBW$54 
@[RPQ>SR\M<J>F,/85NZA!\N0JN@<B[?W1'LGA53HI]@ 
@HRWJ36,T,22/_.GN9:(O%RC%-^DPLI*Z+GU/D8K?JF0 
@]W[#<6B8".W^]LO^+YDY3?MQ'K*;RI!4IQ6RAQ*\I\< 
@R+#EVHK&(WD$S5R75J'2VO VC\*=^3"Q]CXQ0]-ECW\ 
@7ZU4R4(;(]RD(69L>^=CY:T7VL7YS!A)VR$'X!V]Q5H 
@0]Y JG8[$EB$5QBTQ+)-(6Q\1/)-^"]_!CK4_3A;X3< 
@+)N-HQ7MQ]R@J6YD([OXA8*ZBX?5(LU+U\VZI/C]48( 
@=L\:_-.H5T$%=P06B%S?N8.-\^O*M^6JBYOK)K,6G/H 
@D%@.VHQ.#YD&7[.PLR 6H;4,L' \& P2]BHSG$/ W00 
@1IOCB-_X/(<S"[T96L>7/NO6.LZT?@JFM&EKY8(@*'< 
@M#F!CBQ?C,!2>RWQ'%O)?;O8=6(;D"1>;'0)@Z]%MH( 
@GWRBU<\69$L%S:(A=AG9$]1\Z"02GFZZA;QE7RE?*JX 
@M4&+\:F?L%PU88W8&+U9CCSR>FOCSB7*I=Q>.&@ O+\ 
@];VY?#0DQ;'DGCW.@@&\J;]MGC9]-W(IEU3P*\G%F1  
@4H[(3*TY(/&-*L^Q6Y"1VQL+!P6$ S+^0G,8'CT\ZK, 
@5$WT +2M_Z4TMGADB^*ZKD8TW+14(KJ)]2D^H9;"D'$ 
@T]8.WK638)\$$Z=.*JE,-&EN-6YY<J][N%I) X5MMY, 
@NAL_PSZ-2)B669QORS<+M.8%?B!6F<([E4W2\L&Z ID 
@ !1W^4)%/ >Q\3_F3SL/$4D^*HQ(SKZ\V<5_*D4^XP@ 
@2=F[H[L,&[L6UCU:(:\<XX:!Z=(HBQ5@N-X:,>*;C;$ 
@/I2C.1#8$M0=^UGR&B*/$:&\JM"6<Z[] 5?P0Q<IM14 
@<$P2 SJ>IO_<CI$;)RGY0$]KG\488J_YY;+<1>7;MF8 
@B%52$8%%3:/FE<W!+%P6X -W4GVHWYB<:EC&5JEC[-8 
@DRYU&W6#Q4E<H4LIB6G2#'>+P1^T?5S0L7F!QGKLCP0 
@B^CJS\(2+GB\REK+5LILM6Z]XXAEBA-H7#D<E](DN\0 
@V?Y>"A13"A.99ZA!O+. NVG)!5JW![)-7*)5=7DZ)MP 
@7^RLZV;I#:Q&(CN8R2#G"$ +'HXL69S U,T'O'XO*_P 
@# #7E*';0]F<X(T(Q+#W322'7/$4;B,]="9F(XQD0-0 
@R19-J_7[(+VB2 \U!MZ(_.L*4['V)P51JRGTPUQ51C\ 
@*QEF?6121?T$%]#+2MKN+*E$04KG8-:!AY<A4)B,TH  
@K4QTVO,SBFF,/W2BJQ%,F>).<]EJ:CM5#C(S^B6\0I, 
@W)H"59,KHVO+NM6OF_6K+_G%L^#-BY9ASI\/I-#B\9  
@+*>MWF)0V\>9&_9_"E;.X'A(?WUAI(6[.-+<^]0-IFD 
@APB,#D6YOB;C>Q$[!C :-7>?)IAFH*&KF7VM C%SS-8 
@@CK[\!:S4\Y8086H=J7T?>NQ\-8QDJLK8T[!9A)G<]8 
@%(,F8< K.L"MW1<<V!4M.!@3AU@3>;!GW/7R%\T-I:H 
@CV)<Q 3+\+GJ1L*Z"%!9Q4]EQZM+5H-7I G_8Y24=YT 
@I68D#-$CU'5[\[Q,S+/ ^>;;;K8>YHBB*Z'XC@((2*< 
@1W)/*5B((^R A4])"VD??FREC:LX7/@P ?('R.0N/8, 
@EQ']!5K,VH_Y!N&1[ A^+:?4[NL+@AF:<>5X_O[N*!$ 
@HU4^1N/T4^K:]'/*T8HNK._ZVA;$$Q+X]+U@7*RMW9  
@JG;W'4*$H(U3W+V1_W*KK8D8/=+: $D9NPL-/J/'-DD 
@*>&V$]$!40L0MPAMC-(!"-(^:+EIM9?1W- 3;:G-"98 
@;S[/F(J76KZS)Y;$'M%[L$Q3I<X%H:ECG_UD8C&CK7T 
@T9*DF4Y:Q&V['H!T@/:94;1FAD7G1Z4'=  ,A=PU-L$ 
@ZZW*6D3DRTQ<<BES7B,H#;?/IZ0P(,BLJWD)DV[ V90 
@8TH.B0<B+Y[#NM27SYCNX1XVR:+JIH-;C=0E'N)65(( 
@BE,TM7HB3[\@[6'FLSNXQO2';98B.!#M+$VA1G"UDL$ 
@KUB\T4$0Q<(#<H'8D%B[;;#I:.(JL8W/U[5UX YR(.0 
@$>S"-'%!^="M+4A6&1*1JX_4<'NSE8=V2Z>VR8HT260 
@7(=PB3MW>GUT^@,VM3G[1X7I5!A[O7OU:)[CLCP6GB  
0>/H::59QZ;"N3+2&=N!4,   
`pragma protect end_protected
