// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:46 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
mz86spakGytRvWj2O0LIAshn6wXaOqTmihSA8FzfLl4jEPayw/jD5tvk1cp1alnm
1J6Ivxz5PzG5JY0zBXpzUMU7lAJ4fY4cdpKJHGwTUvhJbqHCA5fTz5WHiUXTC6ml
kG3C+Gk0ejoDHvaUFMfJLySg/WRZHA1aTaFa/8Odgas=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 16896)
s/lGb46rX0cuwZl/VuiR4BMV+0DcogckXG2qa2XCj13v6VcHybADrP8XuH0X4Ukf
QfiR7/eMxQPC18i2Kkhf4U/4TQqw/K9lwuPhB1bxGoRs4OVqlhPKjM58k3mjZrwh
0eFgE4bUB8zUxA3j9EYNANHVS9bg0XukZkltZ45AXE5WddajryUeW7H67ApN423u
xxAjiK4iIzEk1BKgtz2Ju3pzx90hu3ZMPjyV5iYHBaaElQIzB1JfXjMeRtt5dByo
R/eiT4VkTxQa4J6jBNPIYMy3txp+V2Izs9XHx6mysu3njgEyJUbMnL/eXdnXspLE
ii8K1pM+jC5khhyR59SmoQu7GIdpCyPGn5thoXVYF9J3e+tgYLRFlUuWCHRo9aQR
tdYwgZOSz+KKUtd+NGZWRY5WpOjNyBsP4u+uD6+LBnNYUCOAb80P17ayrVB3pIO/
T/MmpNqZWVyCMyJo/Uhe7bJFMrl/8l37jgIEY6m+q0QiQs7jYI+CoxwskL2FdHN/
re2nEvekHWZcWPwzkM+MlNbtm6YH0cE0P9bMIeM0ThgUPZQiCMxb+cGSrPaDGZQG
6eRREgqCaeIqLpiEUhRC7SkJaQeHY4sRRgcp2jjpDOxQgR0wgJ65xiG7qdDXMJt+
N6+PRKpvCBtDo+obhfJNTFjW7x4+10f32o5VMpsQUxVWwKe+0rcdFHFwyg5O2zcC
9iEjoF11lPfsOQst+JJ4i/8pxKw8es+QrKkrMyj4/4Y4Q8ID6JG6SYZCk99GzdfO
2t5U7bqth59BjQ3N+pC91tEWCCy9ZjIdJu6J5aOLXvkLw5Tgnn/ONOL1b1Ned0zi
gK8NZKCmqif6r8IvKQe1OeYUACLMT0vhzhtK5ZxIhBGPBH3sp730DMfyfw1iquwI
lqqGD8VD8dsebQEsDxZghxUzDojdCa0Ddr+aaChRdZHXhe0gbTodJix0qdSHcQ0j
ecRivv8HjP8yc4QTg5Jy1WU1QCVrFkRU+6fPfucmWmP2UgwSqL8piBnPxODv1yJa
84lwyJcyqJVLYmNNC6+B/dl6MTla59iani/WFNESYS7q25xP+2ibiZ9yt4f+C+OH
5B2Ziq7YutK2NeYIIoe9A7Jm+dJS8NvBJOI4gis8aTMFt87+2tLPBdmB+deBwNPw
4n/S1n5dN1CHh99ZUJTVhFO85kuaGR0Pw15E/9XjlodG+i0UvkCtqLWBJOkx5wVk
c8pO5AfDJiagOJC26k4qoQ9Tij1lP5O5nOxRTwvtD9NChX4NxbWuEcmmB/zHXnNY
oTZDLShD1ZHUCdYS6BTroAcG3sMSfp5svA/AIW8BK61Us8TPoZhHFAmGyP1fG5yi
R2WaRnKfIjN0nbvD6q4sj+V5wLrhzptN831KimMyYNL/wxghhw1+nzx9H7xlDJB8
L05x17S8NekcM4DN0IOKzhA+T0pE8asaIXzKw3Amif1cKlpGlPx1Ct0JU/uMX3Tq
t1BK385W5rufq+4TfI6T2HdgRrHL4DuVf8bXmKFmSZWn5g1e6yBsLYTfikhGQepH
RlAvy9SxKqSg4Uxb/rK+QLsR0K8pW2nVmNjfSWwDgFij1F9Q6D7LjThJMwjgLgkm
maSXJof3ubUN7itMdYKLsYzdA7tmSeQoPpTtTrB73k/cqkJtDuejEGynOynGYbE3
8DcpyBWm7YEkneKZM1Hy7eZNCSuOnc3KXZSJ59W23ckL4oIpmm8627sJM+DKvksQ
NqBn0pUrPCc8saM9zcEqbRbECi3ec+wEnAZf0dPikx7Umo/4QLB4xvwqM+cKdcNl
eSCOZvRq+bgxFPFhHDg7NuKFmPepBtHEnZGNsz6+7G+28/EAXD6s/TrCr2iydrsB
hr1c1I3UsH5+B6c2RVz3vxdLuye81uhigCLmUVq5kMYxJQZJ18yU2wtFqd+o+YMf
aLTXMJac5VQbLpDDHJdgC5441RA0XPL4ESQfiPV8z5Y1djDmG7smuHXn4O+ZzQ3t
ZtDtRo/NigujZZ/x7c6VP6eDTkf74eavy2V3xs2p84ak0LYLOTNmbOufSm8MGDFO
gH8YVqeXZOhLQYd56ANOlrLbxih5vqu//mfRsN13wgisGuHW7hYWn0QwT+Vkwv6H
1+E9MJOBzrihaOHNuziCP7SjPuzxRxFxK/A7e71MgXxmuLVhrT416TVFPvwPwK2M
2lX+epWPpRQOTsd4IIvZZwn0XB3nDYia+I1CeWWrQR6SOflf2FrJ3YCX90EHnSq1
Ige43QCXHkKeVJBs/hkG7dTnSU239/Mvhsv1+YS2QriX7odByKblnguUzB9ZbCX2
a43F5gSuS0AnvqlXLv42to0eUm8viH6hpALQuUP23Pk0llLoree4zZd7oSwfp929
rOMgxQQSreYlLoSmzYlnveNgzsPmwVBb36dF21GcopPkfm6DaIW/B8/A7titOIq/
KWVDjhpneiEsPipSEqAsr9iKDdijNvV+wBoXviwzBpzhMhGVUMGds+Cs9oqhw/JR
GEVC3d+X5FSOSGSipLSBHUE8z/0/XlPtoefFupl8upkdkmt7+xA5WYYVtrGvY4qA
usVuTabUGSTNSpTzDuSCpHgJ8fUnTnE4l21DF07EjunJRVUudJ9UM85WvoPwunjf
FEOI8r+pWSHynquF9f0do6njuSvQu7MzqQLkIy6le27vRhGbz+NSgM+INwfMB0xe
Uzb4FinoDu7gfu6Yq88R+h6j/4/RrGrm54Jx5S2lrBF8bNgl0Ph/ZI+DGSXGsZUV
Ycv84xFNJByfrVXDqXUq3WVxrPzAGj2w78HEOlCRKxPq7ARXM6EA5rS3+r2tIeF+
nBcGcOpG6Ta0Hy2mrBvWWNQa8K6Zf7xLTyZWtsqJMzRVIQVNEK7tjGLVgAVMcqKw
reRWxDQmBJyri5oRB/TnCRiMzV2uKWv0SJ4rcEYpExoRribzRtGUu1n2wzvMOTPz
2h4RIHYJei7irM9qbGCtOlg3ivMDzB3YGSsTYqrg7BbuCC1vASh8ZXtclu1Cf/jA
pPyQDymIH3axEmZ3LE+znviOQSYxCRA2CHCOzVFzWVJE0vBqB++dvtHFGQDfLlqe
527PsNTs6JPh/nu5xpwGKUldaFmsqmjGYTzxbcUdRcsiU+Gjg2PXYRjPMQ3bMUtG
pO34b7/k8Zdc7RpxfaSfoNDIaGbUaJUUGbYrFCgfoRl45XRWMi3J6ZR7xfzYRMy2
tjpjLLCCK8NwELiGHOWilkuzT77yKnJYZyEg0gQZEh/8JB5x2n+hKACTj3u1YzAI
h0nSBEhX/dI1LhToFUbb5qmANF+O6fNz1Y91achLDw4I6TOhvU0CwdZSe+PYdg8h
sHJ0ZI1PuZx5U9m2L+/ia8SY8Nv7FlFJ+PI0KVZ6xB1eVDjihgTHgHKjr+fkPO80
AZZzq5NNeiS45eSuRLxs6jjUQbo5GR8cGks+DCqLab24x3D/7mlFcrOadrqlLOwb
V8lVKh4LOlbBvTXDtK8att3EcPDreeVlAGziBFNKZSexyV+mHEJlXoveo4410Tn1
QWh71xVN3xhjTBNoRTACLkeotF8YJtUf78Aq5+qs6Je1RfZw6tmHYboBZVmI0xj2
fvIUPto7YDlqSWiB0lw0+HXdMXgPcJzUP8+RAwYkZeFyASbnthMQfPgZ/9kV2Gqx
F6plFYV6cKlmFnwk++SVpodYq68SEk/X7pxnqtx5POqJXhp544CW1/OUBV2YK/0Y
QgKlEJkZD7R6yGTfI/tOwSeYJK2x8dMpUpKGSdTMS+CtQOgXLYu4rhVpe+sZg6Lu
vKtuPX9QXYJhXhG1h8MJgTsIbDVEHBRnjkbekHm4sDmTUFe9hMcA9PzKiQcekGcX
yXelHu3wKJYYEurN25ruGuwKjdNiU9UG9wc/8HD1ViHsEcCzdVjxP0c7kO9XNMGI
C3qyq9cGzIgGjDEjLEmiQDt/0EcZbXTiJ3P1HvuA0ULZvz+fMlhMOSe6cZUcAoB3
MlO+sl6ual+7N26TZ9OaAxaGWGJMHQSOz4OJWOPg0Q/RoFV0vVe3rbpXqf6n/14B
avFNyNkiuFZs5z+857HvCANji4Pgzd3/ZXXAE3CpGPaEe0LfSiShkR46mzn3VwUK
qiOfBHe0MJLF2zhFX2AyhdSqM8Ys35y9CU53dxwoY3QT5+r097zoV3vYq+Kvj/JB
JqA1wHjyGqvTuF7/6ad9Ru6wIRKQ2RxlcA30blmleRq/H2mOm2FYM4Hk64XW3rv6
1pYdN3DrdAq0znarhVmbtUTxZ7NISJotoPfI0FsXtKQTB3qXWcgaBU+mX5Txszty
vHIbSjJJR9PU/a24HRmSoY4YAEXc7m8+aC9YziGsm2nrEQoTroNc6lSVH251eRPh
gLFCFfS7GVtB+mK0QxA58e+xwzKn2FPul7EQRxS9scakybiZhR0cUfRCATHkh6h5
eeDHnac2Ilyn7V7QnpAT5XVmy4qqWK9nHzNHL/MI5tdnOV4yISMq/dVLElAGSRAn
/5+AEzZGY54ds0+7c2aFoPBfotTHh78o/uDgHXV+B+RqqoP6wvlAbzdrCybRB1vo
Troa76NyHzsu289vgOXnstJ26rqFcxMjkzUp7Tm/3mdsrYs6bLA+rvPJVdohaKti
e0pfoI2Gy4zKAoBpOTvueS1dtOop3vGf3W30NxLYd8dmC0SxjTtPbMBzdb53mFEI
JA2piF3w/T1gcdN/pFjKdolYEL18bnGz+JWabanYQRC3tTsFuktEVISwCyi5JB5C
KvSs3RFaFJbWBnXpa4HArxcF/BSKMQpRfZWuD+R/42q/U34yZb8L7SYG86DLYe/X
87CN/uz8sZZCuJCQmqLuQnnynH3/h8nXFUjLOqxRP7Mc1CwZH1uDRaXuwTDt4Ysp
r8k09ujH4XKTPlc0z74oVR4Ps1qxw9bgjCgc2fsmdQCvYOdTesUFudk5Hc5Pemis
aoGbsfIB21+Xut8wQDi3uyiWcE2lB11PeQmhz4RQUzJN43vXr89QcHz62i/0zHgN
7Qvs8vbgifu9tm5WoU2M5X61hoCm053WuxXIighEpvt/mshxYKF8eSkmJS87+nsW
Gz8G0gTs7i0Id4pInHmrklD5t/tPIGGxo2pfamqLyE68CHu141RTPSk5FwUh0aly
KPhd3MMCObrXa2Cs5wNnUMMeh3VSWUeCwGKFH5FLN/d5ub0PWp0oazhkWPD3auu1
2zv3J59ULoeOsxrYqJc/NRdKduyQKygQ3z8H8HxfqKgSetcdu+HHgw1T6ABAt19b
KgvqD0LR9kz0ZCmLIxxAF5K/5qUb8x45L7VA65Bsdu4xDcinmjmEcb/ovCKI0Tr3
sgLcsQifETqh4vbGnnSKlhi4T5Rshr+8LDko+GH2YOb64Fj1/08J778lgfS5H9O6
p+t0PmTLpjkMNa0MILclHLbYOWZgunJmfuhkgWaHFT94RygUvLJFHshCDtoYxYQT
LdL6clRAwh4kzSLwiRl3o44QVz2X4p5vYkYw2UYy0Ov918OhbeWPdF7I3VwvsKDo
6/6nzDZ9Ao4z4yi2a71dT2WGiVygKqN5K8FH8zHr23xy271lE4W++3g5l39Wt3k8
d7i19xeZBhvauRZcFpDd28ngJHdFHE+CdrPlSGQZDecZwTHHqXrfDvFJhigKBjEW
TTEwD8J7v6BGXb68nedoR+T+NaP/YtIgJOiZPjYFBrs4us919mADY1EzjLkADHoq
XMOa7y+IvcQpVt+fFOK6Jz6vwr86P7Haps9BgMHCctdA2dq+iXVMuqW1m//m86/B
aC6gdZYlpmxMJEH9qI8Ui4Ic5qrKaIR5p/KaJw2FjvphowiBRwa7xDytMv/6Ip99
npBH02pvW9QH08pNOeBOsUsqV8xY2S1jPp75AbH7t2TufIUwZfzkAuPg6kCFIPSU
6oNSAmYWqBkcMZlz4G5mAnNAD/8BCqOuuVpnW7OdhKL1aiuP6CoCBYdfEcBX/8rX
ibPyoaENvJsdZDIYHWNxWLn2c2Q6dDfB/CYY5J/W1Q3Jl3XICv1ttbSzJswxWyl5
cJwNXtrQ5Ybg4qaDyPiWkIF3Lc1Bc98qJ5xxHmt6PGtNJWXg3inypjsb+GdZvtCW
skZwqM7ugCC/yx+3jx7d10jvC/JV699UMwS87iSVWhffnPGh70xKpp7v2bUNbPLb
Tijl64c+KwOUX1hicHCHB11+SYNj0G66/1MSoor6ZqXuQ2poOepRPMOQCy+jBWsM
0w+R+3sT9ys4M7TzJGX9TPewm6CKZnOVdSQZl2gk+0OkIkOwDbckO6uJk+Kwz2Qh
hcdBEkVBGn1ZPk5yl1KiuKfW6434FV4Q22gkpvkF2ZxrSbgpvP5ZqrGoxKy49UES
29DLX3w7Zzt48PmsmewqXrdIMl+P+z8KPu5KQEsvioSALBwm+50RembRt7COU1fc
xk1W09ahqE6ZZ+JRTj1RIeFEAcimgaCkUTYQoNF3g4tidD++WHUBlx0Na9NjT3Yi
VXRnIw+DRU/Cz53sAQxglBJcRzQqgxo9sqtpkH1bf9mLvZSuTzCwuv1jGpETKV8f
Yks9ydeSALhqs8F6GWCZHRCMR57XWVQW4adP3jHNo0AVQUSkQ0a4iDfuBxx+r6CQ
NhJa7B6pW4b4abeRWcjYAI3WgMna/qe54HQop0v7iJeUaCNDUKskFlUaRnEGPerJ
/nlrfJ32eQMEgfTpoGdFTnd17hyEg7FTV0xfs0o2l7GAgeVzXngB4X3XQzPkiG/u
kYXRge8K/1rpTESMr4MiSfYqFiylBGk1u3yASPuFEpbQMz9qT2L2px0g/6kNzWCI
TCY/uXv3MQE6uf6z5GahDK4r2duYmhRfDP4TE0wqxOmGEaUJcp3hC9jxs5Z477Ic
xiUENK6v2DfGz+a6tVGA4dtJs58mKAHVetewZyH1hCoHUBTCKc5s+9QxiTuEKIKd
GavdEm5Xp9j4/S6MRER9hfuXU6kZfvqieTjevwuGoz64v2jNpYQaSyXacvZBo9gP
cgiAnuhgidzrmLohCfeVzJbDRiYR+yqOLl4ecoBR4CgsVZkMRpr2p8K2cD0o4Gix
qgCdcfEE+czpdQFIC/aSfEFN0zBw8EAUaylCmZ8H5x2luoi79qatL6ZkEuVhhvQf
ol1psgn4H2v16T4YBPNIm1dO3kQRhzh6PG9lMcpRHTTlaYHS5slu7yNuXnUWCRaT
3r54QWOy2gzLsD3Tm/Azs2OkEabzEYdu8fixSSWwCKHya8sE9Kb2SxJN16XWuQa4
sAj5HwoI+rfMhpYaPSeDvo9Ejrf9M6KNBZQDm71soUimEuyZ3JEQlivzaKXSYbbu
lHNruj5UjspmxSBmLejPhGMapOLXHmLurt8WwXc2MjaPGlRULt+GT+db3kf1m+5j
8+NNcw9hxtFGeuOtHzUL+/gihs374Mkrw7/uRA3NUmEIgPoBkQ7gBaK1T3xo6+qT
0Kma4eyRkywZmVj0gAqzPQ9kksUMHj3m10gdPb7YRVbNIVedxC8f1Pt6kiLMioul
yYQcmLHFnSI+3O5989cD/nwTm8DSkCqd3K+Gl4m2D7zYA2tqWTW74ZcHVnLRx/FU
BDwoKP8Xdoe6YsB7uu3OTQxZwpwGSes6maZnhFMxiNZPbZXc9fd8Pq3I/9GzG0Xv
A0EBV30iW7KLPVFzoGF/VnX4eiFPH9enbHtDdwgvhAJuDkehKLxY4dplK6SMm/tQ
rGETtZYQoKWT/MRojhTBShdNgXRa3/n3lLxREmccRTqT2jR2tYkMN9C7sYYzKneY
qIhyHkTFzfSs1oj+8ab9jE91tzfKkntea9/v96OQAmXtfv5PGq19SLNha8aauPZJ
4fzTyTpEBkCTYQGzJUqd+x+RnqFE6fmDS9VvxmOsbo0lSYMmJYgVfqvtKKypCVf6
jQrJezXF7nNFyiRI4XWtU54dfNicFoUfhsROrzUfjhJHfEEfinWVIz51TYg2tlce
aZNC8GFJZ/yY+waj0+Zd193CsUP6fw9Z2vlZKtAUkgsZj+Tr9oWAdvLrGU8xyZwd
CRksBlduK+6K4kuWFg7s0LpmMXl2AHCCzz1ktPKVQ1F1PNQHY8trTWNORB2ZMLTj
1K+kHarENr5treUJ7dNt/cmd0uVD6YI0DwwoWAfwbWqrxv+wOCMkQ+yGn8rK74aK
IztEMO7xZ0ovRbmpGsiYKP8W5gwOtrA9a21QOSTvFrUhlOvhBwzPVAXP0nG0fg9q
PGyBcWaahIaDRlzN29PizMBuJeB2bfsFykzgvDAj24AmZWB5tKNfA/rLneT11Qwu
Y7IlCggaigfjCMrjC0JK0+LeOwStXjn+fYi/s57w4kDzL4yySFXCJK6Xi8RjoczM
sQ36hpHvd/ZFj8Ye40yiuPoicQNd9GpQqWg03OSOCHHm4LGJTh5bYXUChUBdj5sI
IVIK425cVwkAsfCmi8SwUNlux9znq9cGs6zLUENBURWH4JOIV/mzdJILJGDqkvsE
VXHWLs1g7W4VIki0hji0iH31my65d+Me8O7pXviwkguX8dkr+OO4ox7o76BQvdjw
TjLsBeicW4PMoP0wW8uOuVC/BRAOQ9CJ6n6AcqfEoxM0Ido822DhjifmcUhhppfI
ae7tPWJTJ0QTQtTQ7u+U3Q9daB7LYOQ2yYL0QqtRl4M4B1j3OFtQGZkRV0k+hVQB
4iqOt06qPyYV64ySQj5BX7oHYFIcBm0nZEFGyodOm4Glp4Q6U+m+712yrd0D8Q8S
Ms8MNRACzG8XCVWnB9CSMtu+fqHB2IRtwcxzYrEyNGxmFJN01FA2DzPglWmA8AA5
PAzBsgqlp1cBRnwlkDiZ56LBXIX6z3eJYgTdZOBb8xpoe2zp5XSmQuS1MdRn2+J8
tYQ7s3KYCMtlk2IgoSfmfeNuhR9YDEYv10E1D6j9u3GCeLEMVVHR09/ztq3kW3O4
Zq6mrYsqypWrhpxLUcsqaJT8sHDJz/yfST1VjziRTozyqs5RBbFhtRir5RsK49WY
85Jhs9wiDArudK23drQY/SrdMvH+iqQN1fmG/Ifn5BRJ4LJVmb6scY93osJABwdK
FRmCix+vgCYRWRQJaWNb5Gval2S8jStYyYMxrM1NHgVdH4cozPpRLVLI+Z9K2qt2
CO4paaFwDNeiruYsfjnJG3wcYnixslYkcDDeuCE38stxCZxuIwnI8TKHUZMgWxmz
utlGjOWXJhgQo4bta2bS3RTowXPWRpuvb9H1w9PIXxzufn0DwUj+TNQleZ8pHXqr
Lp+Pv/zD4LHNcSXoNmKLPqHUgwxLv/fJTKMcQvjeX1g8lZNo83WH67ccOXHcaB++
Gcr3FChf3tJC2ywNrPVN/SCv+bxdnmFmua/WRSS6KuU7p/As8KCUEutuhN/hIFst
aOaW9tUfeoUsYE4aYtk88wUgjuVDKPbW0BNaelFiUjlf3ROdzO7oen08y/f+jAZ7
lr5xoYl63hXY3SoFzDflUBaoKQnukrCOjWICxgB2zv3/RjXxgrpWVGdi38YlMEdd
Pm+THFjbWEB6gEq5xJs7d5+Kv1iTYzQmJNi620onf40xY8sHqLLJ4BP1uQYvMF6Q
19ssxIdzbWW4S+di3mcmkpolGB+CMD1avTGQ2bupR5u6UoXWa4husec/Bh1Z2T9S
jNKV3/Cu0ES5Oaq4GlLnKMgqmx7FGuvppw5+CtwVTjOadwIaJ5OsEeC05frtLXcW
AOGAlVnVZfKnJo9XMgXm8DSEJP3QDcYy82/I8WBcIyPXWRNf/LFjkZVHfluiFZME
xQjMJk9P2/mCIq9X1WTe2elzhs1SZyj8vq2IzIlPA2iFz7P/V7Ttn/HyiydxU4Iq
Mp4r7VdGVMHF3DUNQVeh1OQBUU2e2yiAtq0rQqAR9ZrR3BDuAsk4+UfE5N570Y5/
xidsEzi7MWMo9vGZbOcCwxKB7X6s1/1l561qckBJXG0AMZqceFCjbdceGeOMHq/9
RWgmQSo5gVSGsY79UMjsTVjt7yLvpFZkEU8YsVxoQ2AWK/f+A8lN7uMjGaEKsT0t
q8lzNUSE1mFK+z2JSSIzpKDLiKlO6gZDzFMIVqF1x0tJGe4wI59GSOhv3S3XWtfA
9dgrg4SLtMjfJkqOBP0aifhJHhjBI5Ll+E9NxHn6h1Ba2oIZYZpet+P4YZKsUHkC
CCvGsxtNKULR6ESUYXmPX+LgRBTSTKxYBkjRMiwx3rmem1TCWs3nNIqqvtzSjFH9
GFHkXbFZ1j2hKJqzPk1L5mA1riOphKH6L7rbXbYBi8Zp2PAw2iGWFj2bBL+l3m5V
181/shS1rXtzOW11x23DSZ2MJs1/NOkeThGtHvcLl74LcxZqE9jalbpoz3dCdTBB
XUdzrHtx9jSlL7JIv6GgUHSonwptV1SRLyXTEvNdBM/uccV7M6DRswFeo0+uKhPG
iPWanviNLBX0ZRP8nEEGIw1KvgAJ5TdRZqq5J6Fe4ordv4o3nljEe3ONp/LA27va
5ti4GmALmxDSXuGGjPS/5/vH4GwKmPHVA5tTuSXNwMQunvQLQCgAEj/43MLhWe2K
7ajycT05RdZ7oZIG9ucmtoNk+Y+UlRwYcH9kl129PP3Km24G98pMIYd+WIy0QZvG
L34+xJ8Ap02wbDaZ3G6V+rt9w6qDvq/zWBFIZlPSz3abLsg/AEu6+ZIdFptBGpeK
kWf6xxKimmrKLH1NuwWu6hIgcKBTQU6d+mSefN6t/lQ3BK1RhW1iYmSJwwdd6xlp
MzgNEj59Pnewsz1I2Et2A3o+3rMi2KHWIEWxJwNg6eZMlwrqIgcluZ9HBryYCzY2
XFB1fOFiB/ol/TaXSTAlLAeb9KlLQK7PT1kycWeLOkyNeohcnOHcgjYWand+z/15
WDUarhyERahyf3PRo7La/2xknjZeauY+jCARjeIFipyBUP6F+K0efveHWBhQLEEZ
gNNqna51poGN3O4nY6KRJ6GTJ5oa18o2WXxrVpeqoi7w8SHbZqx52pikn9pllMmO
PooU85NGVewtYzUdLaB9FCWABUdE4/wq4oI2RwtbiyKlSpOB2dbITTshV/khQeq9
jIjn5T0ciEu6B5y/pKPCZJcRIWWwmGELWpm/Z8SXlbgaWcoQBpn+lj060Ox6x5Cj
dPwfJWT/8FHl8ZGm3Bu5NBYwfmXKZUNpYjL1+WlPK6Jjef3WQusEtB7fzo/OJ4pg
iyPCtEpZy5Nsr3RhaKKpyV+A8RgS6eszlMkPe2Lc7gGvLKa+9tJ2rD5JlJhBf73e
iK/K/U8QyaLjF1VZT471h90MQPk6MbF/b7VfnGWdUOABw/qWmkSDMvf1VI1IM3AT
lbxKxwd9Ybv97LqdjRi288wloDvAwZQbrSqKT3gR9/2mlkisFPkNn1FxufSvn+yc
mJKgDP7MgDJIsyTwkhYyunz5VST0PlkvM6ZfpgUbkvG7YzNVerROyZgvY8VTpbAX
GVyDm73Z2ozqWPEH5082io9pypTkPibRCYv3TTAHuwINvoQKxIbITOOMPaofb44u
nK0USkdOswK3LSnfGnrXgim5YlVmJ8PRUGyQqR74bDybzyIS98De3snSxSHJJr0W
Xc1UKuRhQe9WHCXh20/C5/QdTk0isfVXFgyc3SYqOTpF4j5SXQvDONoPyOKOzZzx
UEohfBpw+TyYc7HHvb3WxbReswelRPGgdkkUGVm6zMacL/BJesQfF5ccoPWV0Lw3
huub3Vyr73RK+O6Go0PjJPnZdH+upCAGYeB26YdPmDe7Lyo0f1njnzmVGviVKTNB
6zxHBGzbLMN2+qJk6ozgGSqBK60xUCd4apSqrQZoQKn5KJtTDkY9BSodtfcR2/XC
0DdaYW9QhuYeP3ZyBjj6QT0yRJXtGh34cYEeTvWiVQNG4ejNOoYyGIGYNxYBllEM
FWRt62cxbvWIazBTRwohV/+JQ3EsGivMqYNUoUs37S98RisBqvzVvZjrGSZ1XLul
ZMFxv0dRa0G9WICKHrmOckkK/XvUwL4MONuEJ0sTfw4O6kapA59sI/puBRrPaNH5
ovFp75Chdz2XRu/gCM5lPN/yKnnlxYt+LCh4mB4bh+h8KjTc68Ey9tPivaato3RO
oHUBGbnhgqQmd1iuuR6h7cr7qszuHX7darJ16MZROaxq3hUixG0BTc4sAvGYqu1t
vqF5yWl+qG+mkPpHlsx94vlpYvnQ2QgUKkGjH8N/0rhbYUIc68tDzpwdUkisvQOd
DwSONWpdZLGmgwPrgX1O0P9CVJu60gM/xB28cvTX2nIK/IFa9hMX4/I6INtYOAtn
TQEAS4YmGUuLU12nCJvew/lxrv1aVnWhpqjdmCvOtOHRZmCIZCyRs36ENN833E8l
rxXu3Mym2r6uIvDF1LQt2LPDbFjUa+nTnAfEtH6shFYN6K5mgkxOzC4Z9/hZDExS
iuzJNZcAqtBskSBTG4xKAAZdvtXfq1oEOhKMiI9PPyZkj7a7dY/gNEZ8y+LZnnLG
nQdzxhaDjqpPpmjYUmIF0hGKid8fq8oMZYOPqNikHwvfyzBNw7KPNLKmufM4zZkd
BFLOFvzXk4J/XRquJnVRfqQAP2qVL8w45/9afkLl/nWlMoKcHr3hEH1Wy23O3783
uqszMLhHIXGgh0nXWivmbSVFJj+pVodfOeTjrP7d2huYr1Z/hy1U5KswaeNNW42T
f2FkDi2mHyTJB+5/eR08PF1B2uztUri+akwQiDSEfczz4zkdEwJt120J1YNRstea
aemwPObGPxlb+MFIiaoHBqUuNfehUT+6tFszL+VOvtcWd5E6ATme67TxNxUA8v2g
TFs1T2EBFoXwCBWKzyqOAXFNB5DnBwvtYppMPNi2SASEo3/wBmoOmqGIzCfZCwnH
VKO0OY3IzwpRuouEKvLGZg9nTw/TQnUEllH1jQp4qSjYNrngITFDzkqkutEQwlVc
F0p8XBwm+GdnTIi2tI/ioSuiCepZTAOiex7ENSh+D81Y5jbGltx5a2HFTGxZKybc
sW6JULk/2t71Xf/ZaTE1NPc12sibTQxFBO8u+puRcdm3WzDUMXIjFtFpaEWwjWXK
dfyxp0NMCOTrYcbeSVS3Qckxnj7ZS6CBPB8U7jcZIZtWMs8s8DEfEUpLxjqS8EZF
fn9dOse8lz/L8zas1/xkkEY8S+92JEwInkdUsD/0SCYlgV1L+rNo7eaM8IZFj9O9
orqkDhq2C7MRmjznCkNH2tzWRivhKHhsJMBQdWWeIaqDzi2fZCGU/458olyC2jGA
5aAVe4CnsyRYr9hiHFwUrxgy++wQSLZbQe98Kt4nsqjZcOtkfvr3GB2pvBCv4kNh
/oKEKEpl6E2gymMnDo15hhkRcEgRlRx6+cMXu9GA6Cw+XN95fgeN97CEk9Ik1bkN
ovuyAcd/0sKkxmjfFApwTACfGgZEdiMY3L6RmmEW9TTwCPvsTmikuyFa4voIxMtO
2MZRO1szB/RgZKKc806+Hp8nKLqg563UpjE6fyowmi6Jp5Csw2Q/PoAMH+BT8eAE
r8ck5bK+cdUAZFZx6oWY3Qycf7y9gxcC3qMV22VaOenmTcM3956B5L5y1QzJiLsx
ua36I97oJLiXY1xf9IRC3geVWRv2S7UCR72Y5zdHsOl3NHA1vX40tahUwEyXokOD
uLq3ARXRh20SDVVM86sotTWdVDdsRcuiQObhDsJ5RI7+Vln2VCBVEqfbyrDoQbBL
js2dqpoQrNZ0jA9qoCRnBIhUJWP1GGWzBY/7X7PmW3XzlUu2eX5YfFRYgrb0OJv+
GKWMDdhs4caSpRpDtTgwk8uExOpI16la9EyI5IiACkBUJlyxBUiiH7A0A1/dasg/
g+AXigsdSqDpAnWpPqQ3c2ijMXn/lZird2bHZJfSUggXtWe2MYWmlBe1IRHdEzg4
eI1s2YoWZZSquWccCbtMar5h9Mgkzyo+vWEMd314ibG3qfUvnRJ/llrAMgwaiIbi
VntkBb7o6hEaFJAWBc+xHuBlgRGRNKEZPbjiIG02GXTKLcL90pL6JWCLWkzkNu86
b92NY7Xn4QmVKBR6dfdgitV4FOkRuKyGbMSSOCKn92l/kVskzZcO/cXUU5WLCYdY
FkqEV46kmW71jFHXXWNmVwQ5EQCUgk6rtS6vDSZ2c1HQ7uDQnTcxWwx/AjZTcYVq
lV/zbSF7m6rvfP2C0BxLbGp6JUTK2exsjWLCwyDoy7EaWQp+hG9gs6zSSu0u4DOn
g3qLzLFkkiKIu8vbzqjFMj6A2cvFe3SJ+yNh7bH+1LXiYl8z3j8/dcwNUVuMFDIu
9HD7t3ozXE1J0VcXMDpczUZ1cvxYO93U8NOPlohQmuPZIsewREeWwaxdyl/2vXrj
zqPIKBD7DFvbU/k2G/uuuAMiGgYOWXqNVca0KiJHrAfuN77Ao70+pm9xCyjUtcqi
TAIy001/BTpGfzQdeOjoLdltx+YNODuyaZ1j3NCvLOLoK7JSmiwVIijW9LqjRzhD
sDFhMtypGnI14SG5GomkJEJOZJFutWqxYOU3AOGCQdHARIW1SbgbVfk4fvb3WB8d
u00U1D3tYPzXbsemGsOKeo4JxJKVonjfof+sYBBUy29XzyjFLGJVgIom7XWjZwRo
/9zGZDqu77bZb6TkXDdoktRIjBTIrwey0yambkZuqOaPggkVHblI4ZGbHYhzDpJf
mbK6kGRUwF0V0JPS6uqpPQ1pW4xe2shV6qU56qOenzZyj67Zm9Mm8D+h1nXMaXA+
wnkb1DCKgvTnKxsExgV6i5NuNke8iY/kU028ENJXEKYlm6Mfc7KgYBlPF8nCI6+q
1sVsGG5Jt2YtCC5TwPAGrkzemqvWE1T+fTlHNm41ZJYL5TN8u/3En7fZyuQOIgG1
d/dk+jq/++0IBwxXcxBt5koAqw5wYCfU9UfBBH51heInX5jK0avQvJZMOzNRbFpc
sFe6A6sETnq/0GVm3lX5SB0Sf9ROsHtGy+M2ozwEH8eF+z1/ak4YTlxsTsSGiJjg
tgFNuhfWZFuQlgSjIuHU66Vn0jW/1kFLu/qTjQHfvVeclbIOzaJkNFqyxWr/F+oS
Y9JVH00bbxTwhAn8WOEnVTxs1d6VYNHPxeV4YVx9fjXYtfsOcH69W9c8D4A3ni9N
hBTMZR9WuE/KDBpWF+1WOcvm+6ECZ9yNQ2xdKWeUDdMOQ9CVwuNmLTGXhBu1GqP7
cNg+bSeOevSy59y5Rp5H2Iw0PPgEwLL6ai6q4CLIV4WJ+74EAYDI8J525+1MgCt0
ns5cCFV7v2/FttcDjIJqsrbhh0rW6wMPUXZL9Ufu0bx97wI8ZzMHqPdds5hOeskp
NVmJqvFBQTHprU21Ta2pbxOVk6BGAMSFy66gntfVAhE+hkh1YjIqbZZjr8702k+o
iSjuhlAC3AXvAfbUPcKjd1aZ1cwpceYGoSeszez2nf6LbXhfCER77wPRmVIE8Fi0
a2grpzwd6m7/cKCueDTNWgGiXNTpH4c3GLILJg317zWfN2tK6DokDJjUVlqo/ut6
xPNRrw+AeiggwVJyrkuJvDbahpktokWkOg5hCg8OjtTbagjJ6l2o9mVE0Rz1hjUS
KAJMT3bIauS2osT9tKUBw0TH9TltZrZemKFrw6mAnb0TEW62UB6PhzY76QcPa2oh
rPnQHi2b1TrFjR90WY4E+WVXx54UlyVHak8dthcHg/xmNorWTb7RvopN0nIJLilO
s/FIfM2AbpdsIMM/PQWbHlKUCg6OMesQy6bGdQTR+MtAuNrCA5BcictMdQNwKhn+
ZN72kcCdnZSC9ZzwaP+WnECXVyJu/D5lJj7h/df4T3HgYd3+VjmMspZ7rvTD6WnC
1N3fCRKwsGiDGU8j2Knk5Jmt3QC93f/Ned7lWLkZQ7PZLkkPDnweNczVnxNrQOsP
NNUBDSV9MVz2idlFtaY97nWD2TdL+cJFQvzjwRt3sejXZlfR9lMdlPSPic6qcfYz
bBYunjts2XAPRZvUVNQOJIAyMYIhyVuMT4a81uI0raU/sREf0N9oKR50rPNt2hQl
GxYHK5yx/NfQx9TH9aTeFwdVKxuceWaF/47QENzBAJEvoTFbvMaBDRRLGYTRx7Pg
Yxe2qpost+NrWwVRnFFEvlMP4Siyc2VVS/9B806G4GSGt0am6dYf4BzWCyFxxkGn
9EUKvKwGjniq+L1NPdJSrEMEQrpTBcPygvNT+HDfxq+uBCx57ncDSGHmKaSzSXFI
BFk+nQQxStvJMZ7PGkCF3ZLhhWzNJTXpwnWMwHJ85SaCc8Nir57m+scygtHqSIsZ
N4ZUZ1PVMEDOpHCBTAge3PpRDQR6ZC6EjNF3p4ShQDlRzV5p/Tlo2DmCoOfQolYL
z+iUucSyc/wBHLT99bGKPZbooXwAFmXP5pqFzt8wSGF+FFD22ZzfddyDp0wTPUdt
LiUdGutkHrUnU1Znf+CR+3Ue8WR4aKrfCB4NJFIWjBIK0ywcx1gK41siigr8MpCa
3/0c+YKJ0/iAe1vlbfLJV9EB2unCc+TnaPztK3PRZRUbRJF/asY1vFc6UVg4ybsM
fP4DqTKa/mKvvl7gXhSCQb8R2Kr+Q3g0IeMe0cDQrivaBVwe1oR0UoVsNz0N9f+2
NWPoIJexKrEuQtThLXj3XJnwmVufhD/A9ff92KHvv8nHh98lobTP1py4wY6fWvP+
LiJ0xXYBd7Oxl9mPQtJyr48f25fG16nYwweqf5hy42h/eaCIF3VE10P76HKIQ2gQ
GFjx4VJi5bcXYjtuLUe97NoEHqFthSzSoRHAnvQsBoYzBAxGnpMYAI8hrx+dYm0d
p3eaXGtKnXbJMzMkwrEQ88W/9eu7dVTraWtEt0MU1GrAxBO9WPLSh+gBeFGgOpJS
xXgp0zhSzkhyQ2GhFjlb0QvlCIEglA+OClF5rjYKjsMCRZYmGWa3e6c1C/pcq/0E
lmmbg4U292Vho6scZszZTdQ/9BE9fxeZUSKBHp98stLD0kSIppbG3PdZKGNK6wLT
CjSeHWEu6aQ37w9zv9fsC866vakANE15qjx2JvkOOHzq21NS5hfFSLcqYc2EvET2
EyAPQNbG+CrxXcVDbqQrAExwih9PrBA704ofyD/L0eSVKqkga6IsnmmVv29SpbZf
T0/iySBk3fCMv1kiYIyHQHCgvT2Pb8TgbO1TiPFfFSgfufG32BJW1yy2U5+tyCvT
qu1b0DvVY12d1p1FZ8rf3OefsBstqmgLmID6NtOC7pT4gbMOadlc/3ekOQa4OF+S
FhOKieN2qZMax6McPeuommAlaIylmaV7pwYNMfyjmkd+2VSlegyr6Xy2V2cdOzcn
9/1p89NpblGkGwTN4E854RJV7jNXxz5VAv9xYYMhV94BvoZ6I0lIE9vaaSzwjFXy
Gc1VjeCAs5K+EvGMmfYaGTss58ElOTXQskaes9RZq4WOrjWFX3GufP1t9kHv+usA
XF8zoObiIMu0PQNzeUjjPQQgOapR8FCrTtMORKtaqD5s+F5QSiaTx9yifJp3iaup
AbaK41Ud6ge3uRi2DRNqhlVz1CDBGLLLDYyp30FZbcV/tOshS3Xy72S+J2HwjgoA
29wo497DjMxY/hEwnDXy2To1KK9IFqJxc/FP0pIFZ9rUrbMf1xqjPez5QiQTAbbr
33zmsEmuRyUBLWEblo02UAgV/l20mIepabILyh96doaD8cBRozV2953K5LP37el5
IHQI9kiLGFHRXiu7NO0rNXcZ5MEdsDui69CiGzzZFY8Vb7hEcnZ4bpSq3D7+EbtX
37PksMz/i25vUCUj2edJmS9VFA/kb3di3bla9k9pR+sqDxX+NodjBARAmlPxKOhC
UqYm3TO4dICp4eY/l0pOHR1uc7BTWHWtXHIDDC/uyYQbWyY0DADuYI8JLy51tEKQ
R/xacGoHy6S6iy/NReRm/UHUlnO+2wrDo19dcp8hoI1Fvlru1C8T/x2wxgadmlEm
k4CeNaYIHDXVnQW2xWPlY7gep5i9vq0e2/iVqXQj11vEH/vg7BROMKWP3Fbb/FOY
vr17YL6B/gRvHpYqEDx+II4aVaSzLoixo7HIfhzXqXlNrBTk0WBMsZIZ8L+uXH6N
WovN96LxYjARikS2wttOMNszEO+CAxxFwQKu49ZPy4g9TfOXh0Ch3F35eIZq1FgG
gEl7vQHA+UuIXKFj2ALLFXF5v8hdITHsxB4CDYRINOkbbi1mXGUwAMizWOnVN/zZ
uqRyj/AsPqfVBMzdVsp1o7t3moVhSzAn7N3fQekOLLatfS2WdpDIICIeNBZOrAW5
0zmarSAM7Hbl8WYuADJ0Hct3Q/MVZYMF940gCGsFvLuoPbcqbMUIUUb2DvFUG6x/
m09s9AR3WPEXjxx89XTz0ymnzBi7WLMYNzzeqfoUrtJbh7YZTDcuylIj0FdcjLbN
Hr8CjVNVvf/y/KtXs5n2TsEXrIfHK0jw/1d/S79sTCCFm0zTjO2ALQdvfo16sAFP
jC57tKXU5n8AUzV2jFkyl5sf819CO4Q1bcCZZZqMBRBoW7Ti5iorHg3hzBCgbbyu
mD4VrIBpOD38FU6CNOhNyVuDsqfT5ZTxd9WxCx/fqvD3sLTte37zBA2d4JDgDYGX
h8LIMbtm+brhbipgQA0fvgbsFP2jZ5iJHuhGQ+np9dhtsSWit1o2E+V0j+pNGnpn
/4yp7hRNBRSDGMLcVBXjYsCWmr1T7TiPXDNPyzO962xGw/IBupMhrtQjXCwLOU0j
qQGmwqqtztlbB0rzzhX9Wc3k0tgQ2vx3HLDC9vUnZ80jwS93kxrYVOTk1Q7BsqbA
qFukS6iLfQFzuu2KH1G17jWvez8dlbUMJf5Sgm0/8mJjqWA/k66id7GIs7AIw8Hs
wk2qH9ntOT/qCVPwpn96iv4MrEsoAYLRabyC7t/oU7zhAwA+zEsUMrPGY9EHD1G9
OIMgICkYMwxUuLnuFIjBf9mAOm61dosvxIIFDdnQBGnv+31PlMYbe5qdx6bPpJXa
vTFAzLu385OPlnLOH0m682uuQmuo1Ug7EDE1gkVlOs6ZkylK2PqrfK9QZk11nTA/
cG0C/CnqDZDl7BPdMvLqAmmJLThGIPh7EIwqUxdYaMDi1g2KZPfFqqP6FNfhza68
qjTRKwVLfdGTn+0m02/+wiKA2AE9aFGGjXgDK+Bnw6fCx8B0sQFKnfPrFJRNDR/L
F7Vv403kyik2AS36JVuFtKvmR/aVfb3EWoHrJFSs1656f1MJRCmKXKu6uj01iUB8
5EvwX2TbdLwJdYi/lkvZOse2g3Hw7Yexj2qDYPODVXU/U7ti1EZoo0avFn4jt0tR
Fplre4YwRhaODe1wi4o7tyJfKdLFS5GGafHse6LsMd9RdJmnaNB/i8Dvv0hsmOF6
0F0ztRIgmqrVsRqWsIulTeBIZLxaUUpZYicFuxuqnVonOttaG41TOdBTu7N3Zqkg
Zyb6EvVjmq+PETqsba2EnNDt1Eit/7aXD6VFuUiRCHCwNjvAwjVYxYTT6c9uyi1d
JasPTiVd2faWfst0j8GfVGplqyXywdK3zWipMBlTK+PvYQAuoCQkKD3Hi3ETaKb9
92miZKqzhcn1dIs5JL7nnni5KnP8NC6n7UkgKquqJFyrgelgO6ZifXU4C8YWlzk+
NM9srz2tWQqq98EWMNtYejnLFv5D1ewF8N+ZHhj7YPZ3A3tkPiHPbwO2rIRnEmHz
s1wRUMxp5k/CJ49oD8LJRB2fBXhKNpGPi58c1TrtmvBbN+XfqXYYFh48RhLosCxP
HsSEi3WrQtRPVE1Ob+Do8V8Ye8LLUxTO26IGlXqxOWcOb1JZzLVLXhPo3+ESbPDy
lM4GcfZyIzgIKU21ZaQ6jX3tjA10S/UX4urk+qbPKpnVUKI2YJF73yxTaubwY4JZ
sDbGXXLOY4+h80FChiPI3SZLoaRtequkDNVLl7uTKvc9tlFHna5dFqd9II+tPmYK
A3nParwiooiTBRSJkpJXbNVuoJ4JdilWk1SLc+oEp7N/edG2VNf1LpBlgMQivNJt
1V/DkAPjYXyaFU7Aod9Bip6BQztlebR0EV/+Mr26hmIBDu9ukKEINWLvejTT8T4M
b7SHV6XQuR9kv25uQfFo2p4SKgt/Sc52sRaz0Td9CWi3nAwPAT8Bnr3kKVf4j4Gp
XcsgA9cZv7s13imV47LB0n3YX2BEc2IwkIuRoJJ4NMgki3cawS7lzv5xbtqnWtfg
PI/9rRyYi50yrSpNdiMIXsEFoBz5CDG/yIM08bX0aXcHVMIiKccO02vtE3Ue6dTq
/M8rawoIuIiYCIxVMzFQJW8FImgiicURa+rgfVYoqQzsPaHZwYzCj3Kj0W3TirWL
Dw01JbIUv6AtL0RIKbi+y/bUx8MIfXsuXsXmoww/klDaxcilt07p6MGb96iae/MK
jLSzUg06U2XCREysPRBG16Hy2r1a3IJk0E+hitNb/Ej/tT56fXPCuY3/NSf8wnep
EwkHfE353HVyNzWVDrfzSfF4tBcEJZ0dZGYqND29EZOkvuHoZA5YtUwQotIoSHrr
fNf+BiL/5HLhbDNgoYk8me2lpMxQ2BIMeLi2DNxdXxl6tfLbRhXhHtRuUdtHSG0U
rBucLKzMxCVHmHKFw0aQZcwk0D9aRKLt6rqY4Q73o570dB5oRY++ukHwVY5ZT+HL
QUezxxD6/8bhmJiCLSCgT/qyd8CYMDWXPwHMgWjF917+rx0IP6sRgRUEt8GlNIQl
hva3QqDh+/17zAedfD8pMRxr1SVhTDpnAfmyFZXJIODmF7nxPOvmAUHEKU+AdKxm
bt8nzz4vo7jN3HZEfCiErM3RcLEeKgMsSNX8/J6bzHQuNSZ6Y/j6YpWHIVqiIccA
hXcMhZJdF7bAWXoRUuLHhTM/uviv2S3L6GRj0C2K1jrlW5XldH399zTH6rZPxTdP
8b8AWd1jxDHg55ptQNqIwfrNtAgLp59mw3rODQKT3g6zLPef4Kip8pOvACpFE9Ry
7iKDzGkQEq4+jG5Z9xtiEfkBZ9kzNLMJRTmcbdrxuXRBfDeEEXTGSOdgsZE1QJsa
Tx6F0YxcHXmSJEb+YYQpgaYjHhQzKei6F53/niq+vqibI2TTFBTVD2bez663RdFJ
eSR6fi2N3xbuwp3H8nztm2ATA+sTI7Ia5e9U3BJ0CzmzwzgFPxRPGE2OPmsJ7urL
3yZOSt0TvBxMI5ML0qpfdoKSLV7oXaRmadB6tFAoD/PU+ooLZnuM93W06R8Ukj9O
7enw9Fr71vTDUhsNyvYFqLSoYyzOV3IgUvQU73DR4EYMqG33zKSa9Exx9IpjjWEL
2yUs+axX7LKPh0s/PyYWRIcW/hNnDUagfJKjiRrKdNItMzYFiFaIFw1BLy6c452m
aluI9PY82C9g3vqul/1ZziMyJhvf/+2Ikc8RkNvU35pxTsAHJ1tNszHP2dDF+ngO
1hVJFPUpkHbUnejiDFmIdzdtKzKEFp2+fCIwm75co6cnN7BBKiM+0FNheFDBjSAe
BkBrFDUD4/WFDsv9WxelJwUU22RBv5bk1jnWNFIgNYBiCuvnw1V6i2o708tUV8uY
qvR40XmdofbjTfrkoyyCaqH6oQl6C7X0S2hQWi+udbWhpIPH0unMZ25SRtBf/yAo
JK5gam44zRtBGpi+UxGCWHsIhTDzUQIJz42RL9l5BT1274n+0S6HlZmscm2391ik
e999kyyB7t+FKQb4yAuhYcaY7xBZbGFHbJ9WWgi0nrVmRsUJxdGF5XeDklS3Dxmu
+wteS0sroTN+etj4elj8+R7nKc5d6QESErVJyBEmibz08I9r+S/Y3mjm1ji1Btqa
hINOgHLcx9I6tyZBHlEmRHDE7XeTCqoUhX8Z/vTRQSxXloDVkrqDzRCYG77nfW6d
x1UJFSUuvqf/BqgKAzYOLkj+XZ19Jqf2c8Lyq7PnkDOa89Ce6EqpEppDOXj6nyqX
FqIWSoh/6NvouabwlpwmubOiwG5XcPczCG1I9bIY6JXxZydC8L6baN/FtqS8ud+g
l9EUiakcp3szoI5wcuRGjhcVHPE9bKEyd0TMQvhZosDNhN4HOiH0QANvmj5CehPM
Egs6xBi3FG8XCRlu14c9GxKjVNOf9ZJCgIRsWxS9xaBGJFGgeF3GDe2/AMWCdnNV
A8V9TGk/WzDUE+3O+Yn5fxIzZzHGurgghWtDz+Yn6XMWoMWW2gru8zSKNnsU6PKO
uUlW/Q0/m4dsSGIAqYixCWWYGEayTivAiUs/vI+ImNGiW7hf8jUWoo8D24nPa1Kb
2FagY+3/HYfHHYWKquj4zd7yAc6/4gq+LCHEo3Ffqp+aKaN7HLDw8IyS41hFLCGX
bZIpzy4Xi9zAGbEPC0sH9uA5yqo4DdMqmQbMJYJfcwwmWfkgB+nGJoUliGGmQffO
64oUjzgPGCz59ce8CMXD6p9F1Btcocn3rqqZOFgpVg3rNEeGkoADJ19qcBbXIwe7
EWgcaKfTt9dkUWimh/lc6b4iAGymsMnWHxIN2VSWL4Mvsek0bC48MenN/t7E6ZUh
qsYKNplsjtaDT8mdGGh/jqaazRWcedQ2aGV+HXR/x9ZXJquyezIyuYjRFX9qvit1
6cjC8Qc4abK+m026q6oj/QoCZo23o2ESTKLAX394h0ZHjIkQPAx5tf1RjeEdh/bP
`pragma protect end_protected
