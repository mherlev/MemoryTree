// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:52 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
TOEc2CDzFc+JwVhIfIUoMes9FpyRyEYc7foRDPv62cdlpND1H7/AJYtJiJ5vXLYT
STxLFLf9VsnLpepHxyDSMwkgeP8NkkgTsGm+D0fZG0KiFG+aq5apkhng5mrqWAPJ
I/OTxmN/rXHQOB4O740KEk2E2MDdO+J7dTTHfYP3vzM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4496)
CUALyJveSGXqd7ZddhhLYKqPoWvYdN/6n8Y6uVzGanQeidKApIm5U8mbVz7OOb1t
5v73dt1h7ONzCbbfXqy99wGKjeqzEusv4Hm04wsb2BD7CW/4LjjZ0x0g0UuMPI84
USip9y5gkTGgcnru+B9v/WanBWRb8ia9sU70lPfORoMA1Mfw0YjkYMGym4x20Zj2
i89lhprKWdF7zsntsbHtlLv5l6NqDyqZ4zPVa1XB9RJ64ZvFEtjIUnlaFmOxYGjg
DC/eO63TAB1Ibisg6hSWM0eIyoLmQhkOqavRAUrJ0UTDMdmsdYznZawUNtLyET3M
XckzTq44rAnPpdm2r2h+NuDKRJMRyi339YOEPFXzEHZPB3QnNqxBVQiti3VOlr0G
60YKASVCfXtV/jKjCipOQLymIIja4DfVLwvkDND5UBtRnbRzXJv123j+9/tZ0vXU
emVlfT7DecReD8AgeqMnaz4SI7jIddgXxqviRurEc0g4V3rRBoUG4Brd/iKAGp6q
MVET5o29p2ynKnukd1WzHKvT4EupESNPaM4hrOAJdom+W0LhkxdfoKC2aWH8Ka8y
yXifHMutD+OtPv3LJ+56SBn8+yHXPGipAxs2JZQQKJ64vp+TkGCM0/oXlM4i16dZ
fzrSR3Kl5WiG0bUELX7ntg9QmqDQHQR6o+ejizsbfOoaiMeen3BTX49rsXBEE5AC
aCL3VDRxdNdASXSJgJxX2y4ozSNDPWWOiYw3fDMzDXnW/D23gTUEmRgau5rmAtIn
3o0AFSQR0jhllzeWjFkLe+21XZESWuAyJQVQuJ+KO9huv72zJ1tbUJP/9rDHcing
5B4pNixqilVw/JFR3zfaIQSYG59eSYSc92eEIHXYgPDbaOW9mPgUNu3nWna8JORx
7c8QDHnsPksOoLnnZle/zVHtDuOEF6XC9ce0hSh3pm8RCk0OiDDPIRjKQP8isP9w
MLNGckXbZW014WUImGwJnphboVbtEm5MIKRlEiu/YlEKD2M8D3JT2U5fWWOAeYFi
Sne5Ih3MXqjAT8Wclz5q/UFnIUrur6e16e5z7I/W9Lb9bqwSMO/1GRnsI6dw5T/F
NjIWhiXkiKkiKbHWLQRu+hmKEWJuOZGviFLuLUpYJbC6xPizk+AsytPrzO83+6RQ
5DoSBpQhnbpXAVyoyaOpjw2WPjgGhlCG/Nqp1cP0nt+O/GQx4neNQRk5s4MFcTB1
7t7e+WRpXpQn+9FoQ2WPcfADUnCsVkhaD2+EZi4TotBAYpoYwjKs8gRXa089ouQo
um5287vCNynR79BaCZrRWAItFK4yiX/RlZzT4gD7P3WIGrmbYqNRjZpoyGL/+W53
JMHcpAAmmYbD0NC6ABqomogtLbjcCNAgYHNnFiUVoomr7fvBWPOs+nrFVUcFXyZB
AX2OV91zoq22u71pBo9NMx21hXzh9TZY5oSk1tGS2YfqKyUm1QuqZrJi2b0O1pQ9
P947MZEwTt5URJu/ThG89V2xB9NJPOvag87VP87Cq1KzYBdQrQEYk31a4dtEaxZ8
HfU+uCdjm94oD60wQrj7KxzHBu396Uvp7N7unh2oYykt4/bOEKkUWO9r9XUGBsew
YGqsOKECUZOjj/IwNP1CyLil2Ms2jzroyCB0XDiRSAIbDXSg9w9ffldqcCJbmKfz
NrA+TxQzfoyVIOX4NCcUQn6SqdVP8r4obuw50N3Z2reX7EpKfXrgk8UU08Pkovgo
Vnw7IbIk4z8cHc6YaJic5N5X+E3S7qyIuRds+Smh9WPG6iMRzFchuxcu2V7O6+GL
DuonPyMxTpIiq1z61VFKS+Le0G0DPLSb4K7X5vH4lgpY1lS4NhRP4dvlUOtU/jh9
t/ZGdQOp5U0sdIIgmGspUZjgAsXh+62Rkp4etJ9uO/cJnfNPQ5iwOPgBGvvqpW7P
cKw328e0oRZaYQeR39f3JMNeK/ol14bm4sAvHKoSR953F+YYHsphh4cS81rhKlJw
LNJtasgpcGRMgWqmDDC3kCoEgavTcGsSkWE91o3R45P93o4S5nZ207PbRbYhOGZT
Z5OEAIl4fbxW/uk8vxFFcF01G7+oCHe/MDd3qhKc9md7+j5cw3IbUlNEd3lTQz3E
pVzjR/7EBZjH8pxHavYbHYcuXNlcDzrvJkEooD9XH2GgQ/IFn6Xqt32XGO4fsDrK
oOqVQQeaYZFWrlYh58JNeP9Qn0q09XRs0csXx8yXBS0TtzDqUyYGGW7aNqgW6n7b
bU0wysydQqKca2DZyAzA2pOWvo+L5Sdu/kyyr+6RL/0EEeSxWWMFYgnZGoN9VvdH
guuEN+/05RXR5uUMECmQaKfz2R1ENZit8T+JqFPSCO0dYAgF1MaB77PBVdnmGRb8
UweJwoDw7/D5mkc6RabDS+knHQOVumg0gOPQbmkEjmz9TfmnFXgbtvQOQ+eKXwcr
ozzWzqyMHqsjKfv0kk/OhypWOZL7YsBPVFaCoqrJZgagBRus9kYtRcf6cuOayKsN
+LR8NktvbEjN8mSfktDqwpHk/cAEv5JAhYWoy0GFAPBEcki8HkXzsUuoBYaQHPZi
d2z7Bvzm4tdc3EXq/s/zlNbk8JuUVwnSdmO4XKyOdlFxpKru4gaOQeJI2caGsDgk
BpMryrBN3oQNMZH+ESMqFMybW9Svm3ha8XGSaFlR+vGvhWulQD8d+89g2Q7bRgWz
6nKB9IG+WahUVblC8VgoBNDmfUuXLmPhd+gBJUlIsbvsOARSdm34pFkEoZKe2V5p
z/onV9pkqSqIimfw8Z0LGmKYLaKmF1VgM5/MK7WuYCSDR4v58CBOl1vDxNNeK1XM
1CpSKPhAJTsRrl5Qno2ik2mVKhZQJ54IIdqCnZnLt7gHi5/n4875mY2PL4dQYHeU
J6eWR6ABqizpvKOgx1DEyKO79JiNPemjoLgpCfhuAVijbis+aN0kQVppqGNjW+tf
l9ZMcCcveEM+H3UhmNIMfgqi5cQ+5DUHyuc3c7bLcBjkPV0kCO7YEBfl1Vn9d9eU
cHWgg0rMdh8T06NT7T4DANBUExLiQ9UQFussI87nnOTxDAmZYkn3sOTiP4ioAFGo
FkWBBsstnOSRXeN5cHvjROks8aNJBdwsVJ7tkYQD7dDyfNmpmCZwfJffYJBfH3Hq
kX2zjFQBoGCZ40n7S9vjR/TFlWqLwbg6sV+LX+kn959TaTIgsDgzpoXY6F3YFzmc
j+2j+y6J97xQDr/6ZlRTdFZ/1YA9p/KOPjn7aLK7kJB8mU8ODjekp1V9VXo1hton
aD3/UUxjbt/H9/5Y/tX5+0IDlDByz66L01YAv7TIzXlmwt29DMl5H5cL/3JC2ETc
NnRJiRXOLWiPDHe9jc6umN8s4s7dWEFI1DNiifKdDccbNXlnV1o5+FpA1W0Ykz9O
03QgKcWxeNlow+B19q5py0KgJ70sVWBCk9WjGDUjxqR5AXBtaippxsK3PUXzkJu/
/fSF7zxmCK1dDB0021eV3A12QimloD1Tq8acNMSSMlpCBaLND7Kpx00m11NG0SOl
pZCnIZpe9WRqgYTfwO3SJr6emFhmQ2gmfto/M9/pidTe8A6y0UVbtb5FEKQnN2tY
bXiUNMPZRcY9IN62ETAJ07tauoqAW6rW5YBtq/5cDc5cmzCUmJoIY0p67/hk9RhD
fQ1AojW6Mz6zQ+OJLd+gW0fNPOgPFwAsvK0QatebZ1+vuBGdvaFGn9DmMPnr66Vz
xz244+rYsKAs7Tr9oWdWvrcE3UA3m9BCIodoESVJTQlfacB6YB7aTRgsNi1GdpY+
SbsqeQ4HiFsG9iUjfE5eN8GowatRG8OP5uR49AqCYUdulosscKnmVtKmphdgWP+W
7xFIFd9dY90EeCc+9iTZqnBYVlvQgCElo01VXI29iL4lPXixEwi0DNdBD6FRda2u
oN5fzY4vZPMhpAsxKXm3r9qgMxuQoZgp+8byO95xjIPTBFEF0aVtcEJMEchrdhAT
gHjaH58waJkmhFERUiGL0eRIpMrIYtdlz5N87iVZG0w3A+r4f6Ry3Si4q2316tV3
4FW/fo5qEFEpqzOpGCqFSF/KGPG+vcTNXY9+AeGGsT3K2Iy14+0HbeKyXMi45i/b
oEclW+8/gBqLw7aO/kspzYCR19yifTtfM1RAgVUfoPClpjWGbSf9qEmxEqiIl3AD
KwwiJMcBBO+lOAnzdEYU/IMInQ8uZuevtZeHhND1zFuHjFZE7BN+AUuDsVRKZ2g/
R+DDZ9t6423TLVUFR81fncEShots7TyWr+zko4/skOQtJhlbfZMhdb3W72x2+j1K
01/l0YMWJ5kwSxDAJ2Ra1PYCLrJN+mC0AJbu038nDRoLnhbXNEow1hKj+yhu7NP+
AWlWKXIQORx6vFd93g3VmVBblJxhGNRcGW4nGsvvFzT6Rer9b9aeXAccxa3/VSC5
j/E/aRI+mJMy0h2dgl9/5IHBf6NnAKZdMSuTJusN0ZkzW7nWQBHT3NckAeC8M+oZ
Y+7kjK0u+icUeP/+LGRrtqfe5902C+0FzGzKgXUJNQ8ppONtn6Hj3KPy+e+fuiaG
WH0Wi9yHUlNcdCkSPLF39s0FMOohMpdBAz+M+cHnbjQh91vBLubtNIMiA/vKWkeC
Xv1ypsPG0YqhSgfGr6BAjCf5NaLdI5WTC1kPKnDAS2mwKR/xIS08CMeeHZwcqZD/
stC/xmRoDOQjiNn5GvVUo8B1YgpgJWuw4SFcMtUhbPJkdloRB9aAQw9Z68MmCoFM
99ntAA67eJbsZWLhOKZVukTLdqWmzohJv+jZpj6CJ7jmBeAZPnu4thCEkCIbGkpz
3PuEoUTb/urcV/T9GSQGQSeQRdppHgaHduevfAiQu4ajQW5Ia6OW0jSuG2U9ItNx
p05yvFa2SCqmhNwhv97j6FpczWdcpZvbksHFn1ebIDvB5qlbU1pRYPBobk9Czqg2
vwy/evd9kK5mMxfBrwRTjaPHAqho6bPLh5OF8Gj9Q2jlAHP7MS3TbyPYq/NmnB53
OT1KDfDu3lGF4paI350hQVpbT5spIBlGp94jv0P1D8b8yN0v/GO0JeZYwRZiBEBM
s5RZnvr6OtOn5lV0eyhfqtJcilTgKz/q0b/S9Kugef8BrVx1YU0wxrB30YDfVL+q
6jvB9Vq3tbdKFwNVCsgk8GVNhK7t/kLPF8ijH3DVwXfkfSanxF/toz5cZzkgVAOn
2sCtho9nNO1cZfegAzx8qypGJddEzKY/j0mVDd39oOE5xfKUDbL1yjpM/Xy3gtoC
DhSZ35nQSZo7GGc2RcKPxh+7YMXUDT7Oho98rcL9/oPK4HczQYfMvbfZEAeaaPF8
e6XAi5pg/fpFP9zbSzhqhedKOH8Onij1YQJV0o8j/2L5ZWMoIuvNWC6nO12RDZhB
7GumKvoqQHgV1L0Avx5AsB/iSrJ/GjZZN6++uF28vgC5oOBUkb/I2EHapXWRd1as
Fb/eXRhYXru1rLockXjXSruNRCdUAshYA2SnVRKLNDsyxI430CpzS2t3rmoS8Jnc
NEUF5zrZjOoFhMDqdwBDEWiVP5SKLNA/ACC4bO7GCr3ftG4T5dbjVQqKEDfVCvs1
hLQ654Xghw4ccTI0Mq+WVcibTOtj0GpJ95s7dT2r3hLQKt+wYBp5CsGFfke5SPDl
4HsOxAlWH21CY1XeM2ZGaXv0x3kXeXva+pIT79GKLCg/aw+55fkaTBH0acgOkwr7
g2N7tcHvvNJ1eiRyzspNsJ0A0Nm9/DRa5fjxMtroBrYVOgDBpNcnWD7QRWFm0QlI
0Z/IUtyu/8jyNHVyxLdgosDv8vgNHWzrorZfV8mQkoqlLeihG9fpts4XXELRDGxT
v9RWp5hX4QkCQ5qpTrlMJqrGQg+EDFlKmHeMvHnGbCT+VRUcXDibQ7i+l6yUFTpr
EV8T9729F+udKWpQyi0sKyGsyTofhQaZ2T93A101IDeKsPL6kZcINFb7+qLM1g8t
xOj0MnYCkv8V02/4NAsUvp+37qcM1/LNtMIFBJlQHU0=
`pragma protect end_protected
