// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:54 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
L78kLChFvZ9oReVaYSR4Gjsk8n6F/3ZASnoM707JVe2o2TB+2rS3IDIy/gZrGyjV
UM4SDW2Nf7K+shen3/R1o0DLDsVunSvXcA6LPnX1spR2OnnxBUtlssWebJHyQGsb
latGst00m1tHRIgvEXBpKE1AlOJorMQqEk4qmoInP2E=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 47504)
+mcx5avh4zLhERcmL6AAoLerZ17T+pKNIztD720Zt5CmVYEbe3elLTDw69DNeWBD
uc+5uIU2b+08akU3pLA/lT7zxLOnxjYmjqaezkJjMrIKUDv8LFm9SVW9MaS4TJ33
6+z4P/ikcSOyxjcu0fEHosldUgHTbcIWFFPRqFYuf66eS+RwLqFfXpjlHXv3Y5y3
dvqqW1jSZVbRM420Z5EYeItaCItPq7w3RjIEZmrnx1hwRg/X9AA7FKZoGFaTXX1W
oKIYkdm7EQYh87/Eyt5Br68mnHY48aLTEyzezfo+Zx4s6N7M+DSnmX84WqmXlTIc
5fcmH5WK8I1G9KQyruY17tD4p0iI2JDb9NUxpN5HBSKCt76a16GKJLhGeJ9svWLH
N59sKH9W9LQh2tL9GdiHuEufO8b8RuY1ctQHfcs3FjJpRWRUqVcNi8OKQzvGr2J6
slP9uR5AENP1eYbaeXWRQHxUNbrmcF/l1POzgeEWwWATslg8l13LB5dJ8UWdkdCr
ne2tXUSfIPeVx/PH52wTwV+WYq9S3efj1RwTAkgu/FZ2Ny8do4Vrogh1MOmu1J82
xVpbREbX+N/gBi6dkDKxUCUlJxTrTcXbDCdFWuiVDBZ8GSUvjSNX1eNGlaKjxCoM
Wrw/p411XoGSvanX9BayfCVZYqmbxHLSyqhTa+J7xwAIdMmDlaDdcInLTX2KxSnd
l0qU4hRrjnTuDwOowBZJrKK8BSYaCMK+/z8dJ+shSurW4ny1sOFi0Am0zvIiU6ev
nrtoiGXwfvFYqTl9wV26/F3G+eb2FmPaoJFaU5KRJl1CPsuDkWo+Ac27Y9TheR2z
XpQPKHBsYhiMRT0GwMnmzlyTP+UDQRUkLxf3q5sorESisCpQuvoHz+r5MZlA9HFM
e2xSMFLP+LK0OXlxdnBk5qzci07qpAo7e51MN8LT0JrIIIva9QYiUW/B5aE32ScA
Gg86eVN9LmXfHB0jbFHNwPGRd53Qmoyaww3szdyAAeWCdlUYcpH9KV34FQZmkNyR
g0VPd4ngs6MozkHAM3T8SYsySKJSwXw9cW2u4x9uX7hojajZGBn3dNYXA01QrFKU
XZ2v7XVgMClEvymTfwPbYRmowkuK0Z1jfiE3URuFZAR77MOlOhMSJxBElDf6AbZp
W6w/oCw81eeoCtJQGJ9jZVGnLxV383Yrz3KoVTHbP9hgDQr/BuvOOJWIyoSR4L/J
ercmeV24KKmZo4JKi198svLIrq1gthiqrzK/M964Qrn3iDM5gQ3+jkFQDOS2JqVd
Qnh6UxJQinVNgDAOgoKRKETWO0cSRgBL6oKwcjdyXTDzpCY2jSrEkfQAFTzq6Ise
k2jOaJe18TlT6i8dXAo4U1edfGqHKk8v9+kmbx+qY9RJ9oz48erTZKYEeGGNpkUD
Ppps/nqNVpAI2LQEMPrDrSK2CHyGoV+bPn8K1V+ewQLSOMUYhv04njn6hwL1fkn8
I0g90lDyVyYEwud3Wu3Ql7OZPaROTSC3uFtM+bjriA5wfKC3/BxPk+n9Y1Gpfzlk
AMp1EvdF2mg8v8L8FBs8jBJMrN023ojOn595DpSu+pGY40PsJ+ugI8a7U4ueVII8
jq0/lKJWunt0z65AjdoE6HIZK/ZMy3c4bCw4ye6hPaXs4wcfYqHdoGETTRz7kqko
bBKO1szYXHPdxROw3oSw2Zll6LptbJF4/OfN0ED2YE379hpTIdl9RLoFHkHzmqwa
zmEQvqAzAmA4fJdNkSfcp/EJN3qVleh+AywL6DobxobiZJx0LTLYZjaHs34n3RwI
HjWELzTQq8qfipWTIOiH9gndod6N7hBonnID/gCtL7MOcUKlgDE6KC3pXmqvolrQ
WeoPsRDQz5VTQPmSF2C4X4F/HIZACkMW/DUJWWmOh/PT7TiS4K/CNI1gfj5ini7P
LnHizPFMYqRr9L7kpZEyG47j266BVVakVGc1DlWSK5Dku84jaugfxY3GUr/qV0oY
iPIiy9lTMYMZRtpet2RtSkn0QbyN+OJLT6diCcLiGyqkV9CayC2/XZLBdDhszwUD
MqwQaZSFY1X4zAyydwWjwyxwIDIsCpYWOVS6g3KL1ux/tvR9fBOTY6V3E8RW+U+5
r2qvF6Mh/no9qdjgzF1moLyZXkuVbHOc35JL0AlFp9eudg2S4Jond+t0jNZP0B1L
a+vFAKPdfDzK+oKmWyum6+RBdR3GbAkGcsb3lamDpI1QhQOUYBlIdsnINVwJcpe9
5Kksxc62968KV39BiuHirMmjtzGgfH42Xxp/Orxnz/LZAI4suS5rSjOJtD37m2ng
bUnYIf7RlFrZkfHn7KtUUXHosjgAoGUlPn4O7tdWRy3vBV0GKpGefatxDZ6dvZZ4
ptdnw2RUNW5iOv8yB41l2RvOB6307A1a/jg/eAcshmkZ7IzNI0uNa0idE+Dck6p0
0jAHJxTl9ttJiMnhWeJYDzo8uc0ixXWu82QEGEPTxAhomzowWknGq/a4cqEelBRs
t9cXCwHtHYWM+WKu4iQ7DvxKByDnqQEe7oZ8NMe6TtlkPKWWcotky0KSl8gNctSv
GB3rsQBprlIpr87skQc3sca22n3RXm/NDUzn557/24GArITXYf5SqDyjIdqE1VkZ
qIOLZ+Hnu8Y34bk/M/7oII3pl53xHcjXumr4OB3aQWD2uQZD+waGMs1tE03nRkHx
J+qnUtvzo/4I+zxIgxBpU918FQsE2sky+JhkepDsVyHlBbCPtLfsXTIu3spE8ZPR
k6FtdnWmM4U0+qCJjy6mgHlqUZU6/i1Hpxh/VBRWCJ1KJ7VacG4MMLxS99DpVR7A
PO8JQaS6uVYpjjz6nBAH62FRr5AnsooQpjCvsCrGQ/CBB+QuoTV1E+rZ1+RXUTYK
4xJOQ39y4f+05mH3/e85E9u8ucXf29X7a+lFGORbu4uo+Kv4hT7XfEHT96sdlkeh
5Em9ZaF8wG9sbZl3LhF6Oyes16GCLfkExs27rnSseO/grNzOJOw9zxip5kLhfteJ
/R+xPUFNVNkbfXCjg7aoj9lYY3VQriWK2xbKt/cm3x+h6F/F0RAm5mgTMkH13G+K
VG6mDmxfNbqOc5zJWOhETPHNjThKDFhxjpzE3Qmg/m24uUvOsC0pWAha3oQzO+5e
uVJo3rXMnc5ntEtsXhfvEIz+3qXo81ZLLazWZeysXikhqF0OveA3Bjvi3AWnfMTl
FQfkEhzZABrjIaySmJE38ePM3HfIPCjn6FnYkO9cwAG7hLMOM4ZqZjG/rAYM7Dip
EMOl5lrUZmrN8a4/0rkON+1kUkORT5IUnHGwX4Z0SRIoWapmSJb2kf0Sarr6BFL0
AGoO3TMmquDSxR+NvLGF9AHKna5VyvQ/NtCzfVj3sF8mmWGbDlctbL9wAcwczyD7
ip5+INpCB60v1pAm4CPcOCZyespT0FsRS7A9UtDvm2Q4khPMxRs5Wl10VkotOFT+
6u/yz4ddQlki7TlR+R+ypswAOdxbI4RSwaM/cCKDRUkR/ci6u/lZg0EOaTaSqz7m
abCjpIwRc8kPIYiA11MJzRB04599puWmuk9Vzc4QvJWU616wHCFfn5NsnW1+SLS/
0u39uEtt+wwPpDSL/7Xf4Idbrsj7oqn/FWq1JudL9+zUNkic+sXxkrBJilLpS3hA
aUOnRVh4Igebx4gBzeIvH5uzYzrP8Go00j5pl7aUJzBvRa9HyIYKEeA914QZlquE
862XnajAl9d92Jl00h45Ik+9a5NRqTNl0f2ezjxPzkWofUoL+tMUjiUlvAKD2but
1gdRGyeOdI8WUfwmXCkFgoYjxQGNVj9+Kx9wSsLT6HNJ+qVo7Tzx1LRC0RHIEI5g
Uu99Gt051mZbq5WAuLu06Dm8UyjwYyRugsMWkeXxzn5oRDYqDewXyDXZZfZ5s0bB
uO5hLWkwk4+pD0DBduEnjmy7AG9gp3CkWHfDQysBuErhhg6CvkAYsvkwAHfpL+Kv
bYdwUpkJlgz7qa+tjAEE/7+SjkGNuhw81E97OhM+inc3wGptvun4AAWnWnmgbY7C
3Qo2VVfOHjX6AWW1ujKVKOFpEpPFZoIP1QAUEG/hO6JZMWRkM7jHGjGXXrQcJFhx
jfGHtQagSz3k/fCRFnHGUNa1LpOIQcUuzlGCrTU6njfzO7bmfCv4w4GcHd+Gd7c3
DIfCLCzWEihytZ6P5bAivTSR5KIRUdkHRxsqAoNPg++LDlQ71EfoKxLtMIAEUcJD
If9r4LR+iXpnMLLdZH2xPXNFg0Sf/IpTEqjumSwH0gzKUUPAKuUCAr1Bcr+mTry3
+/y6oIgfjy15/R18xjYEAeNN4pzPB1AbhqIYqkKrYGHGzEpKTGWnWgOZ4grBVajm
kK0yrs+xxM+YQj8OY3x9Yl+0LsPHTmbHU0bqsJY+PM6ME93RnlcDZD4ySEMIiK1B
vXc+yTm3c33O+fd1KpmK25DUtUyxA6SC0wPEGFmb6ZS/aOqe2E8WTQFHu8hQ3PSg
9FHTFyx4TVS5nqOFhdmDgCK0T/Il8KMow1NZTeTYmc7CazaOM/SItpY7b3nQIb6E
cbaK7G9xVH0J/1/JEwU0NK78H3wmIV2xT6/OFJV1Yeo52ZK5vMab0iVyRTXcsVzX
fYHb9gZn8O8c+jF16h05FLt3UwGKp34xwzVSq+Qtax7VF/bLUdR+sAuFO0hLxuuj
yOtBESQFu2ebef2rJbZasAQ5Dl6EZeHcu/27AOSoYpEr7JIWGrvtTo1/4mv7rLxF
fUWYUTTkNwEZjByva6JJdpso83L5qmFlmHV3hO+F2WlVTnqVRecJhgZ4eth1y5+b
a7D/P82OohzI+yr61Gaj/ubEHB7cVRfqi6bIzO8D/LuecSnxQtwwTHagjr4IZLVP
Hoa8UmUVOSG2fCWB2cV0MMDCPAQ70rB1uwpeqM3SJkBNuwLvLXnEqdWm0h++DZPe
2vL6T3JmMhcz0oOGWVGYmDIdibOyLYEnnU7yYDmLSekGukFPyylsH8Cx294hndAE
eSJGPYGaBdBxS9EDMWQTLHkst72jzDh1WrU4XN4OAyWWNpUExJna5/TWMsxA5Fnp
GRTzr3sdy4OHtJxp9r5HhQPs/YqCIlr0Imdsua4yvmYf7HWocA3nz94U//L1FcNd
EpemkwKKDnWe0gJTPwECtY27Uy5iQKHy0jsZI5QTkzVGkyEWLoZrTMjXkHcRNU65
lpf1c503mazbXs1X2tPvEW1a61lffuySzrI0tOuP+xlVPTvcddqshlo7hT7b79Z0
B4UrrtxaVPvOQDJwS149LRhOtDhJAYxOrWr+FZC9Za+DooMk8U9tmDsB+flB8bJH
ZH2fSt5MQIVAW1Pv2peFA7N/9OAiI/f4VM61CQhHDeFGyzcxE4UqESPPcjQzGiQg
ULmx2jaLjYKQi1fwKMjuihiTPdBe8MjXW58pNH0LAT9IcwCejHEvVUldBDqZrZbR
2ugRBYd6A4tDZLJvRCeqHMMnkCggDgaD7EAH+9yb5U6ZRZnR3/INdF42iCvXKLSJ
Y6IpF+2WhE14mTmVMURwvUk4PRIJET82TBChERogMkV0l9M0BUPtK0IQuYIYvPnr
AvHT/EthqmC2FBQ2fD4CeOvvG6S96i9a4m5wDYQD1rDEckr21m78mpb0CS3lw2os
kNlMNu3v+gz+elV2J3TPaNl5YaVEWI9GZvtedzyK0px1qDa7IxycDehvpZGlrXHG
YrcnKdQA5xbZeobX0/n28zXZKiefxOBhlftnRpp+s+fsnfQ4Tvc1shLlx7lSdRlc
bSc7IdftefTSGr3idEXrGgxJrvTG5N8gqNHqZlayDeROQd6AvNZlDomrB2Sa+0b8
KS4vv8G2BhjNYZtr+XKVaiPVPING21nN75BPx+ISlNK6iLRrEQJwjLNHQsIPZIrF
rWuOK5pNacS92hdErw8xfB9CfNBA+GkWlD/rr4OLAa1IzL9+rl6SfEsLFuOu2CKa
+AGE72hc++PA/wSngJWdoj9BGldwEXsgVmy49gUktMnF6Rv62LEyrCZ6wE7mQnZX
fPLhZwxtTUs++znlCCycsBIlQek+4UIhwUznUGYGl5m4ttz1FfWbxOE2wRMyxn5m
netGxhjBgAQyrcfOeKCOWj+qosfVbTxU1iinmAjMqeo8xnrieyHMtSOTeujX/BMJ
6p17evdl6yjSKfNFfKETOqBaTYCzEvX5Ac9i/pF865H4ijJdu3Xi9E3cBOQ/VdZq
b5c+V7KPC2LeH4ivKygYL1GJ9R7D284oi2c69dW4kPVWDceuR0k5UuAVjKBSDkxO
Mz1joaOaDpVhopQHCCYDGK7D1fhyRgK2izVNn2WnEM71lt5z2fVb5XRFWsAMigNq
MOwLcVz2h1zAB3sVTnpGrwTbpjylJPUhdTs+jP0f4Vh8L+yG4Ng/t11em//6sNgK
GMa+UpHSiXRciayCO+tQ51KAwu0q28yXivLFaZdVeNTP+lPjDi2zQ+fKblXK4tXJ
/PDhqF4G50HtuVysGCPZ3GQiRi/3Xd8bNWYetQg5oAFy4ILdI7PYEJ10G36yccAh
8ipvfLVGaUC2Z+CaAbt5V19VugGKzxpLj9aRB/GTnrldBrnUe1VYiJG0r3WGkoWA
3VIH5SNLrFWSmF98k5nVJV1QDZMOaNoKkbj/tdJSpJS3wWO5kifsfdbYEUMvBHwi
sNqXCOJocgVcLyfBX26N/cyQ8WdSVGGj4PnT7jOW90sObbgtCO8lOeVBBLGIi8UH
9qbC8Pc4IvFc2gXWsTCmwkjvBRKrU8xwKnn5LfQWlt9yIYKyYz9QdU5NvjLIwFHC
mUHgckEg3KMeaOrLdgSjH0hRKWjH0VEkOF+075yMd05KscFxspYMquuCEfl66qB6
x4akPCOPGCQoVaTOEtsPiPcjOH+VMUOot+8Ffw/DhAGgytXqElZUFioiLRXFAqby
LLI7gb9k8xj3CtFfAqU8zZAx9g1S7DF43OpsoFw6txJoHhsHDg/xJeH0asQwQOKm
u/e/d7Nu+SswfMLo8CxQbckzz/uBj+wjX9O0XubtiNQsUJcG3UorZ8nYBRfRyBBV
daYE0qtuidMkkpYZTIz5zsxRNVeIg8LdHIGZ5sybGE8/3YhlOzocADtylbaFZnAK
URXj+JK2RhmATZ5kTnXtDRVfOegvyEukqr/eTl1P7JsOm/TF7hI1yD26yAiC+MOS
bR2/JKqcU6R05nU5lNukA5ifXzFIytlE68+04OOVhXihz4MhbcOS3nfnti1KTGi5
yurYEgzvVYlwO7kXpFM0aaEp7USiqxotXgEihW9Xl9KNQ1FU0r0mtvFtF4RuTwDP
Heizb1Q9+BvNbjMSRGGjzWnzkpRNX+7WRxrK59x747vzduASjXyHiL4wNfJ1Lm1Z
h92obmLZ4OfbnAOFyvjz8vcLS78vswlzGiYKKtiUhHTU4n2VYA6H8Ws2FD9JS8IN
wyvvPDtUQopFNx9ND9WDVzwAOlgsgqURXF6Ncs8wtfecfjIA5xf5nAi7q4EHu4cS
58R1UaWJNglv0gdhW4EHNSfo4YUQYJzQzisgnvJiiRd385jhgT5H3pN6PFxcv3aG
Dpvz5Bgb5FDjD0LPjqkmKFS9jlfAlPY6l6GY3Q9w6XjCdUJnWxXAEb9VUNvdzz/Z
uqB8+1p3IIW8wwscFDFpK+VGHKUc8lre9saAwJP9Wa3vjPYSHn+ngTrVO7sigtkz
wXUG7IcGj/KOulQhB4wR1XGDWvzZiOAlsiS0JxdUqDXbNYn7KXfTvMsF9dwTgpEE
FQlE16jWnjTSoQRxfp7fuxNHmrzs/40m1wbQlv28T3pAuINk2Z8Gx9qNK4oyoxhm
ngKZKmwaaymp3VyAw8rZvgJJyNp03C0l7xah6P1+MqTUsb3QxPGLIlBfhHIJCdGC
0ftZ0ry8ao5iQsi+crw4/+gzdBNELwYKYG3FSdDVMvxdh3Rp7RZcHRu4BY3aMJi5
KfFTiEi+bYzddr+3+Mtf0TO2mC1x9NWTabRxSQRqg7KTxcLa0rUXMEwZqdi7u5cV
Vz9VBGKz2q2hZ0lu1v9Dgl7lc0i3iHAzDTEKqMccfSGj2hxyPCR+FfhPS/KJ0leS
Kh5trcaYOHcVvJq3B4jYtGsOmSRe71+mLsWG77IYFlFCDqKsMQ4orWQrbd1TLzSj
GswmyPUBy9rlXYpFUaoZ3YckstrCXw7cj+CLCXiIgm7RB3Gve1xVC1VSAO4Ca13G
asFAJ+ZPS7QtGPzy+75222Rlh5rmA6UU2Z6knOy2ltqKr6tBdy07SyueR3LdPQmC
ltkyiQEMLiMxD335ooN7JaU+Sys+1ZWpIW/ilRaE87TKCoAiSyfQaw2J0dGYDgXQ
UNNaD1D0ebO6Fxv3D0/GzUACNJIXdb1hDGDiF8x5tChP0AmqZHI8Dj7bCj2252hK
cCO5pbmHY/9VGGB6Tv/ItWsZOesw3O1cUqprNfOjtPBPwjTRdDMNeC8J81TXzDJE
VWxePwOzY8M1BnAndq2lBKMhQ8dnpkfKBLxNWFpi6NyfHN5Ev69HrKRx0J0puQDe
wwmeHt7GdmQRgIhsBxwZIvoeRSl6UhWYrquWCWaGCgL+vSwPOyJ1FlFNvaKZEzNo
6VySn7SUoNnxjPAWocf+y/zAjtUX3rVHQpNpLGtypfxRGpWrTsUKfuM0q9t7ACsY
06NQmLVuz1dDmi+mwJ5V5OD2vvJ+Oq7ravrQg9autVOjIj4e6GmqYs9MfSjl9wJH
+ROvNPQPCCrigl5JIxg0T3pVkUzm95r6rpvPGCrCK9zhFJnqoGfeAAlBdUswf9yW
2sgmrFRHZaQq2c36zRDIifdhYyONVI9TS5tXM0raoCCFDE5tPqDrbvVZAIOHL9Nk
OJHij7HP7fSsxrbxDytgArHwlL90idWJGB5F/mAx1nGXcSeTv35xKeAg4Cb0ayU2
RHowurALapydmOIf6xX+J9MSRJh89EpBD47LHxm51Tarx9AgExSDP8+UT/+Y/FSy
dY+bXY4R1q7VffZ1KWLaSNpdEh8ykj+ZMnLpo0eWq0sKbzDiKLFAv+ldsn717EyN
vFbw6mQBjQoXEp/9LAC5N9Z6j9xfFUH3OWd6IoL+gu4lEqc1X11U3X0nAMK32Yo3
JaXDYy3sVp3n/Ic+7Il1iULA5Q9Ieduvy2jkfMR//HsVfm9BO0IUolFk9D+ZIgTE
VJfO7KTglL1d+biM/xfIIAPbyXooFuOzn+0bWmJKGytAZiB710BSGQXoIni/dcU9
O9wUh5aOW9QaqKlVFm7oBmKVZYBxwnyZUrkX2FxpTe78hgOH/Me9AwRicrPcTycm
uv7aDlYRQX0EuBaFMHYqHqatXDMLDkjtXbVkUhPBNPlkD3h5H6Km22xiUTZLjwet
aaRFQmqAJF8mrTksOn+dgybF0Kmywua7p94BztrVwIRnHOFphc1uMMwdMh++uh+G
5lXpzZnw4taiMKmjXUIdOlbA1TNx0bk6biHQh2haNC0t6ll1qhwGxcYbMfwOv3LA
AORjjvDyd5qoQcFcllNqQbzLHSrwbGpRNT2IVymoPnNbJKTFnRPT2Nc6S98mVEhN
nSgen77Biha6s8aPBVRNMX9Vqoff2la81JKtQV36gr3C+J9WOw7HG0Y4baTaax+8
wpiU7yelWp/PavaZ/6G85ifoZMnMxOUnTvCLq9YKkMDtXbop7G9DNFWNwlvwXlem
oB7VCiMxV33w0xy7U1aRDjC9aYHRxugUSyvKmGaA3Y5PKC4aF+xiY3Yd1SqxF4wA
UZ5q2mdXMUx1Ba+37zMJl02VzWbzbL24A8SAZ4NwCWOGzUgkgZqK90Ui49erEodT
rZGgnCtMCGjD0qV8VduETTea06RHGQxGcxu9OrI6SQLdqxY6zgysJD/vKFozvc7x
EimDwcfrZe8n9v/MtfrPhcN80XroNF3mdVaLsKaE0flpjp4rAOYY/EtxnWDKZC2V
zjoEeDzB6avHDj2zotkjhi46tQfmFhX3BxEhgyeW5B3prUz39iAj4DMB1QG3g8Y4
KG1Uk5Cc8Qx2oNwdTnPBTsFrwXFmiggGac9ZqZfw6esE8D7R2gabEHyzcFqyVMYb
/6jWXLTBkihzyFHekfNIp7mNItWRr2wv+fHPGRE3iP9MzWAT1jwRLtGAipzAMdg7
zgBuWLDU1USvUMuwS0RAieEcdvMxrqkrRFJ5Lxh10M4bfFV9qNiquJEEy7EqgJSD
QF2X5oG+Sf0fVwrT7i96U+pveOyeRyplX0C8mzn6Tnm3c5NrpdoKNuoWSsuSV/SL
kU0Gx1o9mewzcUb/lQZsKNavro+LXQu2ORvI6ssrm9FUe0jOi2HRsY5D98xXOemG
qx+ONeGgINvQcb+7RNwd/TxqMENfIuEXT22JNBrJKRok1FvAFVFCFYCsN/r6S21C
1FLOK59Q+X4lB923W37aSi19WkcqQWLTE16V7rLjdU8VzTzjI/Mk13P6R7NQBrh+
ZvdROqTljXOZDLkfyOFbVT51G4ppOAmytehgoRGLbc4zsROVjE3RUVwko4FDrVF/
PEJZ712gO/TSme8Xzd7C3jvzBE8dHnbfl4YoqFP6WjxBtpQxTScOLNOernmYd6Q5
KOO0eQ95XcxIMzLHuej6QZPb5Sk1OqvvOIzJWwxXCA0qFpGr0L6+KzooNus3q6U9
hKMfvKf4sy363Zrp4iYNpjIACBMEWzbqLSRdUdmwQtKv8tGEsRxsnqJqBIXeaTbi
DjVFZ6+FFqpdm0EMOEJ2TP9LNU1nSF2+7qoNlS3Tk9F74DbKZqGjThA5WAml18+V
zMVqDa2rre9BhnZbBpAudNvMqFESos3SfxM2C+v/jkrcXHqydEvWg2U53Tbd3OKv
cgvAcMJFuGWRCr1mwQj0iu/QGhkOwg0U4djEcuxCgvMwVmAl3/y9pt8oqtNF9thg
9Cz0p2RmITXIyhUT50ePYv0iUeX/xQIbvrVJYNDOxxhspeX89wl27MvRk65NrGHr
8zWwUAUx1WHVd7HZ8OWaVu1Pkpc8ljFJc7gX2VuuUHOp9uLQr8uEA10NXMl+PY6K
bGlecJFkLhBVSp0Vdeg1C2CzCOEHPnxvxwyInOPOpXX/yIASYdQcf4sSPYTjGN9y
uO6kNMSqP3dW8Erh4WzuaRrfMYUI0hIm+KFQC8q0EjzbvAJQHXHLoQLNrAaYcHtZ
b/dQgGwJ+7P4OFKxvZXQ1s1iC4lgdLGXkpMwnk6UiPWXjKCKXiLxVvQ/jJ+1uhme
zQKpJcSdWGmjXh//q/FFKD7YkLcCEJDJ+b2RiaQYLpRi7Tpf1wNMS76+fWgWU7nc
YeYudrN0ytZHqbeW5XAQ9OFZSKACtg/4rp8ICwwMksvZTYLOOM/oZtaiWaifjQ2y
0A5FbWF7Wmf5oDgdvoarucSikWl+UNGxCCeAyoJgWNaQAAX1X2lSMagLfsOGvXmS
6TOMx6iBsT/yiptxDDPuobSjzVtnAtCxNFEVfdiUqAys0VvgdCVdPadhOHKKrXeQ
b+dCLbfey/XujC1VKoIYSZjz936GyMDDfR3bnUAIt/hsewCtpNubUtCyROXjmDjW
rhCQsbR/gHYqw0hPvfnDtc4u4AX7QHzua9bg0L/AHsG7sPQ8B1R9/qBLoCOWyLI9
fHE1m1MwtlVyoGe6AqJnV/WcDpAO7MXADhSHbhmdki+K7xcH+kklyV6w55H/Zb7+
BQo/XJmASj2hAMQ4Vx4I46vG2FQSvPcBERkiYbfXFUp8k/MRWCf/ilUKawWZ0GtF
w/lmzY4MBt6Usk6IvuHZXlib4CvLGO9lgrubD9IvGBB7NMuBthjfe4Lv9PJ1GCKr
zZa9BF67Wxp4IA/V4QeCNsm4tu7b+6HVEc6kpb0n1WUhU43MKPdU0pv3ciGWTtW9
+uRNmsY8bdYfjmvgwwHA6vyD9Zu5mcnexxnJ0Z0YMfdoW/JIU+xFie15QWjITWsu
MBgEjtq9tWfU8VP/tvrs5yzvBimwjaEYi2kGwJWT2c5iC+xn0ULZdjX+qAcz7qDm
2Vd4Q9v76rwOtuTHtO+epoVmn0I7Rl6rRon5yXXb1LHy4CVC/023i5NT2i9MVkyX
Hw4MYbbBc1ctyZWvJMgLUQg0z1ZF1vetqy1G4Sls/5aIxV2QMkyRSfaaRrQwro90
W549SqGWMDSsGbHQn1qT8bKzLE7eT5EJ7SekTdS+1wbyptkKV3q/rrJ/l+f69eqH
FqXP+2nIgE9S4A0+EeuvaaTL/WvvOB4QxRGyPO1lbP2Brvsr/ZMeItUiOqx/EwaR
hsMtth7DBj3GWaH7hJHlWjN3LKusauOLORynOfT0/7qHbr2zpYeez16UZuMvl6O9
6wsQpV08Gg37Mho5nb9vn7kJQpyT5amYNU+/47s01ZLjWfLAUeqCLOAUiiTIUk91
ngXdidN+EB/Xu1R1Lb0QrQjcDntC1B+7N0o5SDzy8W+5JHPM2iLLLaOERqRI3TyF
GKbc2FfcaZNjdmEKF6XsSmqO8OYxxXjsQd6A2DIQrCzFWUoGWBTBZEhP1IcbvD7O
cYZL7npUpu42LusM5nSaPhtlFt3oPmfcuu0Bh+OvxGoEgZZrIM08Jp7E0Ej3thuZ
u6Lg3CtkHZYDK1sUObE2Doi78F1bDvpyhXGXGgWRhlsw3eXw30bHUhFuwIs3da86
eji4LhWj44cR+rh+E+UXTcQa6W+Ozur9Ec7hnbFmGXJl+0fsGrdMsIkh+dwagpCK
uxZun0X3g3hdRfdTsTzaxnwguPkJ4VAjXxUHbW1HByI7TTpO6BFTiOB3MOah86FA
9uss1ZKaAZGH9QiEPcf+2i8+7MV6a7alsm4x/aFOyhadpVTquqpOpjIwzEd1Ph2H
9MrldCDEc/bhHKBADfKXt7uSLR2RxqblJguvsMs4YAEwZa+q3uS3WNXo2so27dm7
oPHluhAZTs1I628XvS5dPjAZNoFXUIixdVxnpXvgkcDSd7FMeYmMhX1yAQI9zWVu
uTzAL+w5doW2CsXOayZzBGtVc/bjzWXZJfDcdwSbMGXZnMfs6UHh1/2TpLjgaQH/
dJR0cQQ++PKreoicSn/y2lVwSFRskmB7VRfL9It6h/FzxWyH3K9oUEaUsF7C7dBP
lnyXjaWwMnmZKgXAJy3Ingx3FTQNxKBMBYnrG/hYRDvXTs+LPldEDQtQEkokXSG+
jKTPL2RxYRP8SXGzmpWKLyu9y4cnQGIMBTZ0veKbuAJvnJKzzKCps3RlBPISVZUR
UMV8HGACtUvW0I+NQKTHfYE1jtLVUlI9X4rPObLnko7tkdQlOAClXAF9CnCBfAEW
KNjSVOt2zlRtkwEXTzaThcZhoO+yn/zeEObOxNNi4YUfmVL+UU6ptnxLEbI2vd/e
vFNUVo4e3LSXqQ5tQv6PpzLceOdS96XAP7EwR20JMqfdJsTBVJvgTVieFAs9f+u4
Keg0/8v0nOdHmwZmZeXPD0vGuV1HT5vR3SgVAP0UrwHLRA9SANqg+O29z8Jq31VO
FjEwNT7/O7uAZamQ0z/ldIXjnfdkZ3LsApnX0YdTBKIFcDIbMu1Agyf4vlCR/wYp
t7ce0oACYLs9KwCO4f/1bfyMLmC+iKz0DQxwzIOHgdDsB4y5BVvE9Oajp0qyiRAQ
8gbK0s3sGIGr8w77qLN2bDeyEhP2iMlzUxO+0esDxFYjF4FznVSSnjdEzQyvmq55
y09jHZHDIfCrqNK7duegKT17gLADWjCdOhOB7P1MMuNMYeFAOixJhZPwZaeVwr5p
ZHVUufwlt71y6xC8OEOfA6Sm3YHFvpoC3w+0OY1PtXJMynSLTjUk7Q2U8eDbd7VL
I5ab7Ib2orHGoMpL9qPn8RCAL7GPtslWqOAA3Ooclkbk4bMcAL4xPFSXigbqvO2O
hbsai7VlNJFg61ruf2B2Q+SgXdAnTBidbtLNkurOuS7FH3ZJM/VkL2ERsGxndhd2
93Rgic97ccRaQPmsBxbboGBIlrzSKck367CedKpwsf0QHWJptHtY3FXAbOlxp5vJ
gNOKcG/80t5o0SdxHFxt05xQdTwyUBHpodRHnmPwq83j+QM9TkG2qoQMs1mzXZ8g
gUucYw13rfKO8JgesJA74jDeyj5xI0z9e2tl6eXy+MCAJQ+LBY/G2aGwn95zyc3S
fTJu72lr8eYCocRtEPLV3E1SbTQsRgw2ZwSr9EXUm9B01KIC9FVqxzygaveGOdED
RXV6JbHnhWAjRhCYO+OeIWood4fQ8uTwzTpSElITEio32KhvxYhWwuH+Jem+H2I1
k21E2JwWziDxYpybsKmwoTlilWLK5rrVmQJQMvmPMhhd5XCBZ6OYJnO4RlFJxNee
huDWaeDW0IZeQ3oRI+hh/bHaNDUj4XXPIurm/3YSF03Idd9JiiCsO/S2Tz2WEnBS
s+MgdsMLWs4xyAf/a6rkVVOrca3FLCy26ITxT63GxY4syEykJRTyLRBMkAU4PFPv
Q7hAl4a06qSH92JVES0lqj1bEujuAfS/I3YqHfIUosQ2p9uqXN4yaEUCP85X+d4B
atqywJtxjI3GUwzGhBuV74CFSH1vFbHYfqnP5SwMRVAjOtddlmExD7LQq7FQmVGi
titgz7sm3IVTDX3TW9m5iJZSE/DpObac8IDyGjH75w93dxRWgmFerJj23PEL3FAN
rRmB6WT5rlZlB+rMX2+ReEZ3Mo/lJPDxva5um2BnQ4AtTRD/b2F1vu0EwNnb1FN8
yk+qP0ESwjb6M4EV1M+MtfX6/yas4UweeWeoLbHB94rSXsTYof6817Mz0sA1hoYx
BRTaIBi3C1+XsbXkXov/diIa/TBVqq9wZMkvygpJLqx2j4G7rGb1b/IKfpMHZTOW
Dt/C2ec7dOSFZyHXF2kWWhg4JcL0S5mmmiRJturEPUIAseZWMorF5lohap0EPAvK
Lm1dxRTJGtWQk+LhGZeHV0YaVf6IfSSQsHIMJmHQgPbrT69fTLY4Ob+/QOfe1Sg2
JZRAVsHNbP0h+WPjOOQJfvtf+NwMlgttpcftmEOHiLVJr+NNWpXbfU9H8c5L+bYX
M1J9VoNCEiKiqUuwdfRuHGjzRPa/UrJGEF3hb3yQB8sh+uX5QwiK22RMtiZ6uf6Q
yz9COhI3XVYZvG2U4eLqvOwlExwDiJPzxF5K3KD5z+L/XD6F1acnpEARjAgNhQ45
C2xyAbfGktAxpWAoXSuEmSd/O1NNCi6GCOcrphu6J+p83XuPFQYl80hFAfxqRW//
utH/jRZSHU0bOhgyvA5C45skUe/B/rICXm4gR4iCrEEnyrYINZDaGr0vxG5KHeFU
ams2bJSGVB9V0Y52KnQyZbyc9Hvl1rf/KUwkFLfw1uY+x6k+RAY0HO2ZNWA6+BtC
tnm9dguAqX+MaMdmP4akqAmoTvmKmZMX9EI/G7iiG+QseLToM5lAomEIB5p6e3EU
QEMfmJm6Bd1lQLNUP9h49xhhqegbKu/GzoRxY2CN6UBh8jyRSyMSMNC98wsGmUP9
K1NapfpDH8XkusnhJXjLoo/MkDcWxkDxOxCwjNG9V/wt6wzArd5rV1CqnkQvlH+s
wNIyaFXZSSZ1VHzf2CQQi8FUagUGqMEu3IMAKLnKbVfQsJHtwF4MisRTFJyK4Wc/
U+TThB6fSCiFz87eTKBHVxSHexwVdCZ4T/VxkseokjRGW5G+PfNUU0r8YQ651E2H
kXYEHz9+Md4vjkYbOa+o1E8XX0qNHdjQMmaMPzZNy/9g0bQ8LygObBvCnsLiz4ts
9q2c2p5kVaOMkmleoLioKB4LeJjQWKFHQgIiFbzosc4elIuHFD+3D/1ykMceO0rS
KU7UfzlL9z4Cw7jcfW+haXpZxmD6Ssqn+vmNRK83fEx4l2xsvw0ZloKfZw1lGOCC
TvJwb9zTkV1wiX96LdZZ3NuBhtq/S5fVVGg3yyLd1uFi954r4YFNzu3Ny1lUwf5w
OD6TaeDOEAAfTKkx/sH39FwBJpQ4AX0nVCTsK2czA5MGjg+EvbCpri0poGW50feF
J2REo5y8lH1pEqAeGRCGDfvsAcbb4+jjppB8iO48C4LvAnLbP6HSBHI/XB8k6j8o
i31vXBs1pQmRa9xhtJZfqM+5cJB39kMnvE8r3mOMBy3xNi+gskG12mV/X7OkOT6t
XolbV7kMNL72EwmYzWuTwS+qvM9aJbzmuirNPd3/MNjoTj5d3MqevpRC5YpgDPte
71I8PeYZJmzwKcfpalyQVMgnpxBj6ov2k0eU9F61mWDmv6dYET3GibpL9dH9JFRY
G4e6chy9eSQgaiPAa9pGAtbTMNMtb+ZG0XZP26qmAC3wJMOsLWfsfaau2uVfsYrO
PS3Y+MyZi+tf5qtslTwMeWTiTsoeQoW74MvhipoD5BXoEzqGZ8RNiYAbJ6IYJ994
aeIXczCp2Ndkp8jJ/Wz9QyZuLm4j19R6EgZ3dAkYGfVK/puckrCuAPKQhvdRuXNL
wDGyvMjH22SAuc5Kj5jVEOY9UAdYpIstmgwrXoUq/FBkIXEMiQT9KjvNTSDkH9+C
/DNZYN/fOuv+DH2V1JLRR6W9ouy9+VcA48++S0v1IoKSeyFp3+E72RBXU1EEpTKq
QnP/toYlrVnJCu3kOjwRCTngTI8i4o2ZAr4licSZTIXEMa2KJYU/wLZcNKleTiEd
hCPIV4FgPogfhAm18p8x4eIfI+ZSKGyjZtkBW+c0u1BUeBG5HmKGEAeVNbCstp22
3tpnpcS1TY8sgzASt97QYmW0y+RL8INqgMgiCqL4X5K2lGQw/XGSzUJ+7pDodAkk
0dX3K6mRR5rdKUdBKnwnvThbR/IQeewNMQfCanKIvtN6R8GvnWzbMRrJyzO9Y0xa
2jDnJyZ1haDXBnXM1ZixrSOyl42hQbsGB0GxwkCUHRdoExomj+V9xxKovhNfHRGw
pN1G/fh9yQPRMF5NU6TGq7J9DaPsI+0YnBvUsG+gYMzeN6x3Abukx6jKC8KX6xCt
9LQXqqQCJ2GneFxbFgEM2ps/dOt1uQDPCF1swdotRv14FX1nHCYlMxjtGa0mAMlS
Z7ZgdmpOiKZEgGrOTkChvVDnPBTCT103yA7irNlQBkO2jd7VK5uqmcEcd5+rnbFH
17Ys7I37qAQDLtnNWwFSuBP8m4639vM7vLbl8cHuuenmPWGDwyE3/BFqkUwa3rDd
F5sdooz84B7kBR4t440KcPEU6SAWs6l7/z8iqeUqmbyAVZTokBNvJDTF2VFKoQDo
q/EToEBiHUrcFBRmMF0Pmi3YU4yIQFA7PLpP1dox2MKqDUI24CJr/mbY+mlCejcZ
zOEobZfJBcvmBVaUeC1Q0H4PZhDhgazQGZzgxKeV4JDk23RmYV7MTd3omVlWr+qB
o7sNHxjozEJ1yMHtmVdSDM+LGPAo6hzLeEDiWgDHzoaLcXVoOC59RUwezmjpkiH5
xZWgVVoEH9dy2sKGyXgqD4ap4Cv8EdfCNojVD3xDGu1BVQGyaqkG5tpearH5zd8B
JxBQR0XOIC25EsCp4EU1pRPPpJDpErD5NdaXOmab3uD0BrljyFxEKV6M1Fut2KkW
6aPn2vF4490AsfXsVzrGv9n6O0ecjrPg8s8CxzYx3kM0WFXCVcfKHUc4c77PTjbW
oymn/M+bUcwEh0f7KsMzKFN/RPSN2szu+ZO0fVRpfXcoj6eUg0AaOssTWScJs756
2TkbLhDoOatdze4gEy/DEWNnijzSSlEsIMJwegsfVe1nZows78rLKLm8cDK5Gyy9
axeikFwafnVr5HyxU4gD0EMJb0xMXvJxTKAGTAHskTIgbEPbW452aKyOfh4Y4fP3
HZ/3s6TMyYJWfcR3JT7wNoCf3xtZaR/0jL0/gC5wUs5cIZT4SBrpTkk0TaKzYUS7
97ENmEG6SeLbA2/60gY8pUQMhc0l+0Qa9edslrEUz1Dwtdfic1eAELLIXPfLf1DT
ZWTRvckBjo/hpFh4n39oB4Wh7D8cKqEtIga0XfgBU3RQJuuc+uV9QVLNnV5+vPVx
T1NSPPMsSbDlaLoxiGz4xSiXd1tdqNahKGzdpZ4lwoFr6lZZ0sN97APYJQcyxwju
uJOcZyykL3wl6x8akkIz4JRpKf4Ok1Csl6caytS1/igKwkJqZt6veVsMGDSZaCu2
NgItrfnjirliK3me6D9AVq8sR/uFuuj1QE0D7ns8HkthBLZvE5IxLDaITCA18ChI
E5GzC1lvt3QWBlimkBsmhvRat2Elt7MloNwMkn9+DiZqqu2bY6wYkMNOneQ2jCfb
L8Jo8RUK3cb9ZOSNAhcIRXIsBG9Qt53xNLJEGrWCWCI1rx7k0JdO7zjC/pM3+Xt7
8roDEb40PVFI/aDRzNlmtFwEX2TDrSlwYHfgnsDU+JGkAVJmJP+TUEYIHVyEwK8e
7HXkRWqiQV0Uzbm4IB6Lw6HPzK/mlg9id/jvmvcTSnBRQnxAm5B2gGHBwfG+teNS
vfd/LJjJzP4RcNsfJX4MQOyWNekVi3xlsrsR0oWS11deB47/LQxOnb6bPOj1e3Fj
cLn1L9UIdWTYQNkD5SXm1jixPcBpyIQsjIsV5TuVyBHgJtn41pzBU60CcS4kN/2d
j3mazbUPiOPdk7Fw2ApHWuKHvQKYgeKW80Mdp6n7Q/KN3w50vqSXPWvKggmmzrYp
LUtXp28Tm9uS5uFTfxyFz3DRdE1eeN+WavxLd8nR+vkqlkKwkVpXWbwTvoSDqt+F
2tL3/Xq9vORRMyYQ7CkmK0qQbV20Ab/aA3ADiD9MLiQjeigZoo0yw3Jd4uOIX47N
dY9rnhn2b2VfkQ6MiYuWna4ah3Qqd4hwjOZmT1wcZk3YSnEbieMhIg+IfoPw5rFb
6IVnxHrSqLAGpOWbJiP4Qv66wFNJeM4TmVp0xz4AjTdJjLaf7UE5ZPt2lzMyFSS7
NE1KM5qLt4SOWW05Q5nZTFRj2t3shoQ4nC2SUkDMQRc2aggxcqOW0fSIF/QC0Pre
CK4HphgamMxclikEjpGsU5FnyCENoXIvopQwOIOqVdvmh08+1QpONErJkEqPFU4G
v80IdAMA6dzKOueP60NB2+YsPtPewSEKAOoG5YlpoeNUfmjX7E+QEd++fDub/C7Y
Mp68H3KscRQPCySVATGMC8NoyqUoqIP4h6sbUn2JEG7HocrDWb9uqop1NveAnUD/
vgiN96erQnd47w/45bHq16dIt14A/SomhdZlfoY9wQaHWma2DuWyrDsvrg95/P9g
Ollt4LWzpR2BFWVcc6HSIUsziwJsKRbnBZZQURXjFCIeyovBPNICHXxU0BGe/qup
Oo1ElRrGSEYy8k8F3MCMwlSPAQFUGuZdGo8razIYsO4eP/wbL3sFlWSg2xaPp9eR
TY0EK6J3ysazL8IYhQBhyXFPar2BQ52HY1upDouWM4y8XGNSokdeSG5U0duQJslv
DfLnAv5BxqTnt6yVjJQjNej+xSbKXsF5mEjev+IzI52G2luOFcZFt6/7pMJNja2O
PbseB6Idu34fhXox7kw5DUX55WXhMrDDD3yk0sv+BGivrYKlWl7Mr6wDLfLk5vh9
mHo2kIXRTrlRVVqpN4INqEgKoeGgZ0A65meney8+eGTKUphjcFHu/8ZsbIrYeH39
m4wlDSDtoNmj5sGS4CHxds1FBCMLxoEUOlYSm+kqfzVKnX270E255yPbDtoFB61M
7BjdGfDlmn5Y9uuw6lmKornGdNx/IgXv3HcXdSRG+MlnDDZd042hFjd3GZh3vFUW
wj/oWC5eHxdRMagUPw8We4We5kFLiWh8DGdfnp1Q9yZl3//M7OklgNu+JQNYYFs9
kdKRqHv4AIjNr+X5DQkbFysKJEtU1R/ZH5jwxLjhKBHqpRK7r4iVvyI9JEAoaOhC
t48qAD+tOZoATF2xtO7AbsXNmfj9fQgC4H/nnZBef3VBKNBbNM7E23ald9TGOiYQ
DNIk7vlIhhfJl4igIKr7KV9mcBz/1lRSVKKW0wK67qElJ7ziYWGuRgUefoIqEkK2
Aad/Un789rVqRrQoLil3l6/1ChGzgpv0RTPo0nh/FIrV/m89+Kah6gkAQATV7mnF
V534rpT+S+zxJqTJkM+o+m2VR+bGlLS6c2f/3VAMAXn+GbyWBjksvZiZc3wR0jMT
pP44cDyKF7VtIHyy6mvZIBqDiEnN/i9E5mrdyn/tnP6jTcByfsL5NwLOCFqrQHsj
I7GKy+MYfsmSCe+7+Lp26JUjUTFkqfqrnfaONWUXSuWSqgf0huIG90zD2cmwytZH
EB1JNg1jsaeiMjJDWe77KrAqmehfkoxE0lfaCKiV8VwPwQnUWlpnpytuFDITx+1W
Tq+6O4IcRpsdVzT/lgB5XO8d5lxE2iAT5kKga0hrjutLaQgCfhlT9QKPcdL9zFSt
FsJCdmqnzFjA80mVKETEtkexYVwM5dkFqS0cIk4VB/UwfH18kHnLDlXjjAcWHD0H
t25optVyvvPUk0K0CRwMKL8O02k5VMPVDxZFivU5Fz2L2xSvQJAFbZenWn+ASDeV
UoivUnVps89npfeAeERHg3mVCN7YjWxynHjo1jhKKXVCoAnM0CoQs9w0z38DQKZq
AaO347yajbSlj/g3uYdlh53PjhXMAGoEBLFtKA85Xgi1GdVLaNnw1gRw20VyL2Gf
2EOuZoUnTUbtwlI3EnTWya0r/SzyZ6+AspCB5cfHdpOsXnjQ0vmUQr+WufWwxMtT
1TfFwbODZKaqqi+J/cUuG+XS6jXJABXxZpxi8w1TIaZs6nnu+JS0/P7W6+Wp7XBf
OhPUJj7z69vZRqtUaSqAOs/2Rp6lCnOnLRe/AUDnJEKKj/NcTzPnvxeJ95W8gErD
eFFYpq6oyI+LMGvyIJZe4+O3+nSfMPmXD5eeu/9xohRkBRfPlRU1aYVoXbMBgsv4
q5rMjBrW45jL8PzZNBxAdYjAq0OKU8AGIbdJcSQzQeivXIXT8FVYjP3fDJ2Y6Ke9
+MkU1kK4DIJuxYci6mm4wUCQ0okIF9ehnOPRX4cph46yweuEipU3w68qABqBKfjr
ZwiahXUxQBb22PlXN3JOL37xflVVpOyNmeid2JCMABZU0c/DYbODAM9kND5odoVa
DpiJjS64sC7Jq5HyTXDxE6JE/Jeg/7A49B7WpwypnZpi8Acbban98+Fv3BJoJD9t
P0F823osRn0+6vz/oU4+Tttjx1yTw0A1eYq8XJaU0eQNj97Cf/ABkCoa/i2mE7vo
R88x307+8TBc4hYsjyVtbJnmlFxT6nLqu10HYtePDr1wcL65CtBltaDwudvseYvK
ZiKkgCkE6VbBzt3LPneeBaL2dlT60emS0zFGLVwsysx37MTQM35xKdVnjK10+j7e
vW2WO51U+8A1hUyerUDATO5oUDFB5/2McDifTROoTbXtQ9nc+UOpF9UKsb4JrUPC
VD3KBxrFM+FFQz159TWO8HiFJischnyJCvx3qHwFhTYymT7WNd1AqtWIvDP1vMd9
XNfYvo10ORNMc7RIecl7p3hiqwlOH/mKmZWTFdXuPSBoJCw7R9ChvGHU7SQRxH2t
LySnTOFm52XDAG/4osXjCqHsiMpJaGdk1nzw09aWUtYQ5ulUv2t5hxIfWYZqSI8Q
r3Mc0an4YnWsIa0nJ/U9v538jcoBPP6LOdSPYLk1laMRHzCkTZ/EwzyJVrUyNlJj
mQ3SM7F2bVMzSiyPfGzB5Gf4xiBTRSUFF9Lrld5IxH1R3zqxBU0oVh/aN+KgphFz
cIazOzrtA3E8gkEOvZhcPtcQYCSosG3ZmiAema/vlIljiALCYlWHml1nhqFWzVXK
v4IZvmKLoEXDJeeF182IRoEJxOIyLZj3D+0ykBve6OdFIhHR3Z3LAQvcvOrPvuJc
qY6QmdURI0rNkq7OiX2ndy/lF1Vnwvw7HIFh3PLgPVNzS8eyHRR3/dbgTSG23KV8
WF5AvInU77mydoOhE9iIkLUv9FZ34wQWg9KOg01Jf5zU+MyGIT69Tij5gvACcXPj
tpyBy2DRxi8XJVulCD9K5iDeN5Jl26r3A7lZ7EP2g1zgksVi8MrQmsulchZrQVrQ
7wl5IGE8rsUXeYKjKI66C/2hjpPtCTc/iQ66vwz+xasQOLmtpHT1fGOW1F01jp5T
CWd+qiw5YFomJ2ShLVQIAlzTBGmNHuDUj66AcQkPeGjUKqNyEzwiubxip0UbbkcC
lsP58x+O+kjmrkG2rh7TbFGKFXZZ1fe0afJIAvYsG4i4jiUNo/lpfl6DTqtQMKte
40aWTiA7ox/Wg0Ps+/w+uc7k8NZDb1rKIdiY4n9dXZlv7SPvymAFCu/1289KHIKw
c8+SuYTyDSBcVNy0SsQMmAhs0afHASaK+ZE4YfXdTpspWZXYJXs93Y+eB5FwVybx
VVPiRik91ukfyiLT4soxaqjnzeNxDJnhyh1DKDyf6HkmKwmuzN2haXY4dl+WeAug
X2oooOxtzhYKDebZnsIGafNwTjhrwk9SlK/XBve6dA5ZMUItVbQY3vqR+PCQ25ZT
v/C/mag55Qo9GoWpTacsqo6qeIm611WR3Fd6DuZt/Ix0Y33cN9ifNFV62wVxhP7t
vwMSIPg2MB0l7KX7cGFWlW6FXxvXo2GT/t8mHBwt495wUpBBJA0MrFg7CpXR0HT0
jaViixC0vU5jwdatJQ7oU8y5Y7mWdy+w2AR0JW0IZ2DmQQZ77ROc8DhOSXPxXTAv
UwWx5bn65clQKeN2C1X1Wzl/spvDc57S63GLN/IoaTxbatJbV+h3qDzZz2+D3TLN
NKkGlTH+sZYXZTyxAdmxIvVu23KQZC8Fh8TCqq8uxIriNLOES4yzRZ2S+diVUX6S
XMCBeTil1k1QM8W5Lgm6YEC8LirB0pq6YcPW5QvIgfWiRA7GUR9C18Wxs0mKr7PO
hu+ox3BB3Xg3GRlXdAsy5OCGO/yRB22/IvKiw9YTYRRWXf9jxxeEfzKsmqlfjzEf
mc3ji/JMREm1ajAFix6tG7O2MJeYUtvo+As9a7eJ7oCyo66nbcI9SgC9IeA8nbcO
igtUdyurterNDIPl20LOlA7akCLTyRyN/htXL6JmFAQzmn3MOHEGEfqlgaVO6ZLR
gAEmDA0yWVh+VwosUx1Q9ngITObtxlzD6hbSqRqcgGhooV4KJnclOVt6GU5ANBlt
XNkIuHHrI7FEdfaHzFAh7LUtsU9nn7gVNomy+TsXZ4ETMM4To3tyxT4iS1C/b0bJ
NB6vmKSDI9/mKsTxHN2PyrNv+WaR3HHN31NOCeErVBu1+7VDBEs0KUoWlw48nAd9
HpGR+HPDJ9MpGS8BsXYQD+lDQrrbaxIAxiuSzAG5NxZAMExdZDKIVY+CS7ZA6Zx+
InKKl6qNrpv9oDGst3U845rNcCgFtogAnmUnGd+dmQSXSd+yiKeo/pSVd15Aa4KX
g6zzmDSZ3TjMGx/aVMcI1DWiNEbsuYVdmiU+44MbFYx2gj+FCYo7YuUHQSTsYjpz
xZe2UNRdhu5K09sQpTnY0p+GGsHxbzMF7QuEbjwbOzAKSTty/1Uje8MboNtMRcY5
IQaoChI7cD4AT25cU1jsO0RNwpVBnBvRNmlpSvF9bwoTrkl7+FsP1Lc3Obm1jFD4
5c2tPEMVu6bgUMMKY4NfByTGem8fyQDqA/vgtR5T7v8Fx4lvQyuJBkSp5H31pMFr
2o8Zjr+AEPwcxJi5znEEFqGbsycoNGj+QtH/Ex/olkalWE+Ji6zcKQ6amXN6t4K8
KbePBhMiH6QWHwLm18cHy9ni/USPGHFc1wuBr4Xz6ESIR827wr5YXAzQh6ijbCuX
RAb8/QdYsFgfBbsErg8UCOzE1053fS8HiaIMrzirC+BrOeoPtxqys6CrT7a1f9P8
R1zwnYJLifOmSpk8EmEZce1R8vwuWHcgaNA0HKcvwTsz5aVwKISfY+1kivqOophM
HETQEKJ6Z2/8QB2MHG9Ws6riTyJ6Q/PpAbJSMAuTVY59r1pfqVQhfqvsOOimsFXT
/AAS6KvvMKnmieyhYhjBkJJdYbCe7jf6MdsrDf/FoCaoM6pEJyhGtskMphTPQcFn
7ijIMMIbecTrimqUxh+fQ4PMe25r6E6fPYAnnFeFdtmmDHGfigGSC1pDsujE1MUf
3rGjLQ02/Ec5vCJK521I658SHrjFL0qGgnKocZa+MRl2Xe7Z0j85XdqPbDTFvBhP
4av31Z2s3rfedNQEX29G9wCfbznj6jhOEWdFS46NiDzT5bBZD0nX1cBcl35ckfXo
wwTHUNH4rOyKD62U5hLtA8LrY8D6Mr7y6Q5GRWclkzvytiG+B0/eGgZM7Vq7rTpe
h5/4B08e2IQcKlLnbsqd8CAx+xnVeBmCbTysWDKJT/lUNUwiaCFNNJ/mNHEVDH2h
SkN1t5i6FKmHOqo5JO1X24punYriCGUTZ56h/CirQr6ovRPyuuK8ufkK7+8VM72p
bHxp5g4LsRJNyMb+TYJrQzS655AEAvOMQZagBOUBmh7WWiGcvFOlTgiLLdsJh8AU
6T3mCh49SphlO6dxH/4wdjB2eO/ZzXIHAXeEhvRDpLCIAS5ra+SnOS8D0tS8L6v4
nMwFdhvIQggRvxtKh++ZyMXo/BGJ9XC8x6T13VSBR3xgC3lXTL5H4g78RISY+es1
7ebvKT0waJEwvm5zpEL/R4riRPaIirVVxk2eNlnkuGSsAYCG+mGvH0VsL6XWY0kZ
pjJZUlkA40JvOvrZOHQQQVOqXgh9fQIt2enC3rQIpat2xP/bv0R4BMlD3oSzha4e
jAspaxXNwG5ICR5i5zcQ10LhDtQfY/Cr+/Xy1RtrJmy+KpmX1eeqf1n3/ozasKJm
1X8Eha2vJ2TQPGMxJcvFiv1YTkQxIehwL3QWxf/jmja4NiWIHgpYTpeDm6vPmA7M
gVXhlTEE/gPhb9btAdkyhTLx04pvCrtv1OP2FvaxttDMHNFpPzPGTE6VPlt5PLFF
VhKwOny796DC6ytgjtGxvpszwO90wVMB0gWWwsmiSMY9G6V12seiwmxtXXb8TxTb
GrDjTD0DJ7ffIvC+9eAi/VcBcztmGpD3RRL8xTeDpaXRtRDQd9urQygKGAnVFF3G
mf752FX7PNJ7qMxTnHW9gzPNB882jI/s17MANgt9ui0Qm+3XPtPUHGDVWOFVNuWh
57MYx6uX1Piqsc/y7RZ+YVoH9oU/iwe3enQwSk0g4eiv0WaiEH/ARcwLryyuFfeZ
hNunAgvLWEbhJP1qeCfrqsWNgBOmeq/djGg1F+72H2bQ3S8oqzwYXVcePSqJHyFE
GKqbPFO9KmyRantVDPR1CmRwQRjoN2IYPhunCC+9kMjawgNmeGDSLelhajNvY2ip
oJc0ZxuvjaX3V8YCsAmLN6KG5EFQXsiQ5biz6al5xA48iKuR234TXbojsPqT4ll2
pEmQaYz+IhDOEGvk3RUtwvaS7UBwqWNnLveSsct+P8vwXwsQ3avvLqZjL9sdDW3U
FrV/lvS/QLbBUzlyyR1LTxtUGoOVCELl7KWeu8+D+t3lRR6sZgTOZqTpFLvGrnbc
VKepNPDVmL+c1cpaZR/9o45hc8iMhWiQ1Q9cp+ldShW/klRxyJe5wAbSi8gxbCAq
aiIfg9Lo+THlX+2z9sD2wowaqdhQCRRdsfhlxfYppwoXyFSSjv7F4a2yZyCF4aYT
LB3gMMtplpuiEdY9+BFWkubnJ3fu+7sUqzGZcPiehI9e+PXixXg9mBmCrxoKEm80
+QlGvuPsMenwvZW5Z7d6lvwBqlOmzgWlcH5iIpHB4fi9/6VvrDPDwhSHNNBjnaww
JXxjhI3bi2ISDUxuwlww5tJRHoPXZLubGU4/Ow9F18HE5zYFqapC0QncURh2sMni
72eAQSDee9K08qJS4i3NZRHZPKR/uICgaTtSmOSkYmjBjwnlS+tiIHINz/mt5IZI
M9TWSYWSyJQpC7KcR6BDW948ZQjYo5TPl7PPpO5AmFIM06xNc96RWT4ATDgNhPZK
qN6QQDja7vzRR9nackMxmZH+//JGVf63iWEnX8Mj92wHk/HrQ30dXDnB0K+Kmqzw
WGTbraMrj+YTdcu2TB/dMOgxOC5O+cae/mNbYtQ9vRxdzUqBaK26pinrqon2ouBq
QhfMKQRfOHin8/q2BuXUc7gn3V1zVetyBYjCSYimeA7mTC3TVGjJlpCt+RkdmZcL
HJC1WzIsOdvNHHdRxe7KgX6ra2GpM09S6QTICIB38G1Y2cmzzAJ444sMtcS78TpL
VD+ohPgLzTzHuM/CFd0+e/GDUChC3uPLamtKGv8XbBDc27UQTsPptQc/7UxmoT4Z
lJsZC2O2RKwod0Ro32dpyJKmGQo5uUhIU8cexwPHfzxYhNpYD//WtNvzbUeLekfu
j+ttyKjwPxMci0t8GPYao+6FzQtURsgyyuCGcc0fzMtN7h3eid82meztvMh6ShRE
WqZWqE/OJyBWCE1ljA9RDdR9WN3Bq0FFxzj2X1PlLVWj4gAyfA5W18DWHFs/NsQM
oIl4vKyZL564hkmZPoQc4//GGQp1+/qu1uSyIfH8TzV4jdWlNKlnErk5mQIaH64A
CaHykeHL71MJfbMPekTwK8r39pAifS8FxF40qKiLDrKhw3t+sNQ5ArohqfZYw4RU
6ws/3MU3l5ZGncS/k0TXoeiZzkQdrmaS9M27mRRU0hMMbg44qVZUL4gPa7mUYtHH
AjuCLQ4wqTrUEiVqD/R4lOws7QotG5P1UdKZEpRMm9nyp/cD8wDVef5x2eyy7uzG
d3flOemPVDd2/5KjQIsqAO08p2nqD73CvsGES+aP2YLegSjvNV55Apf9b3tccB0W
0RbxCmRk6U/5tiueQTwbK/E+AOSrs9KuaZc/3HoDs8nR0LNMqUS/JT8mlkX38hEg
xgV2uZRYnAhj2y0mCnXCkroS/6WC4w6WpnCGZiH3D2V26R36+/ZpdZhGpfIlxrV9
oJlvHhXB6GAmEvvZPg23fcLVn0nXbetdRWJ8Kx/QBaXTFiaJepdMQckLbDpzVlmO
hJq6O47g3rl9HW/eBa61IqUl/NzEm3AmQ6dkcK/AK0i8dtwzpzveWnk2hIRrStEU
0K92IWpBbgzdKZQXtcl7S+37VITGFbvZOz2shaYLZ4tP8BcYWb7mG4cqAfDExQir
reZgpQZ1PEjqI7R4YemkunLypOPmUdLiPQyei0USHJZNCtqFrmE/R1G17YFZKhep
WSkq0HLfL15OUrCi6LK5dEHIHFzQZNlZLHO1s6WU+B6KiWxGEYPgmHOc+8YLm9Aq
h8olS+lIqyNYd09fIRRAC6B+r1okChiavcjjOVgR10G8xElr8KgA9GNG2XVcAvuV
7al70hO79YZecPeM3o1gzvu4ZH3miFXCHcaO7xYyIpquy3dAk3P8DdLlAiPLWNR0
JlarLVPwbfVzAB8ItKXBO3P6JO6Q3tXf+8AJxtb7gJLRvsYAf1gSCnl9qlLz6OZj
asj1O1uj4H76p1EWLMaDm8BLjlV0EhNBAWKIoLvV5V+JFuWQ/3Nco3ARIcbXF31Y
RNARWpFpiFyjtaKPnt2Y5Gz4TxlobL43javD+Z8rAL5y8cRE8DqLb201h89C3mEz
PWYbYIKZGaySyy501uBmp7ttSqgvXIlLkshVxJSH2HkANnFVWVQq0NJkv8zcb4Au
7F932g3sZwSkUntVHIX376aGbf8hkPKhkB2jxk8BzJLLW6Dd8gQZO9MVcoTXxL5I
Co1GpCXfQBbYnghU+2ImbxEK4RLNx8R5Og5lH+TdgK5VPfuxF1BNTaNXPN9WOZsj
ulrDniSZJVwrTHmIcZN/qWzjOui28yi+qMI8z7RHBBgQ0FANYj9vJLoYzwLqgY34
bTDGIxPrGW0jEOv/zBItM5hnjYqM9FmLhQnrtE2TGF8Nahw2/rMOd3vA8/y1iXI1
hz5Af8z9TrnZNMvn4C6C+0kBdx5GzwtC5BITD1ypB0NJ3qFVJJ+tBkeIq3COy7JH
XWFwZPp744gXgSr0vu33hYWa8GVcrXou5oPkLlNCaHeB/JDRMzUR9X9GW5FOvCPj
dQoUvit63Q1pXwuJW2VmvAjwO3RKETs23RlG0RW9y04yRGRp/qc2ej2gH6+xnmVg
c7yoaynHN6axR6uLuyXlOhxbXkSKbq9sEDmZy6OnlF04LZdkuo9ozsMNPR08OdwY
W/5azpqA1XOSyJLY3Zh8Ipj6dqL/aEAz7MoZ+vVcVe4epGtpElrjmFvMxKClWDPj
wCZrtUS31qOMpFiu6ECDZj8uLHkX/VBBtz379CifOsrho4DPeQp735tp7CefvfYp
qCDrdp2UaadL2rLn0RH2DAp/4ks5RIHJtJyL5+kmUmAJx5KW/agm6/xvMxGZuKjU
uHu0cP/U+KnB5CoAKt0Myj2LKwYeC96aGor8cSmiGFPlVZ5//CvS8IlQfWagWPV+
0ULJk025UYh8HfqfRg9ZC3NuLp4K4MnjT8+PYs6swPldsP261y+PqB8HMDA3S+cO
nt0vsa7Gs3idUiaPVN6Lm5LE1mZRl+3/J7F2h8wWPA3dGr+UkwCN39TA4XVSWB5Z
8rGV2hTFgWZMI4nMhtkZWY+V4jTy/PRvoWTuwK6Gx/rVzmZjHBWfovcfY7CaMq3j
e0E+ourNt5BEYXuSH1ucoepJkr4YxPXa4YkFxLe+pJNTHNkYK2nLH8kCPilDn3mT
dc5yJ6OqcNL8E7epByu+uhnXPltsgiRVfa1OJtA9jSaf1xnf6sUYQSEXhAn3eJtr
vnLL/zrOVjvljc10lzws0051pYYtSFznnOk4VDRA5oXb2ZY1YNEeHJIyrBBJz4Ko
F/j8E+32GvjP765xFoznLknLMAc67En2fDB0hVfzcxhLZUJIkM8EhuzdKRkfXp+T
KPtzTW4g6mhvDJsvt1Gz2sXsHxMJxLZZGTwF+ZrbdtznyuyrUZYhKu+eFOh4Ofb/
nPiJR1qUjrZ2z6H9LEEXbPwxnmn9maLFGZTVn06p5HPR+rGcSnJ/38V/unPJVr4y
HZjYmzwkvwxMvecxo7GCWBeDmTYl2mU40cyFoDjVqz6R/xPjGIP5tFHdalP5ZjUO
KqcypZYmRJ410wk8iNMr01FZuq73x18ghiqgzrx0hvkgV9Nu4iOcy0HRVhLv2IkV
wm5i8xdSPSoercyM8lQYV38p/IpxJKYODTee7RQMRIJb602c4QroWZy0bMTzd4P/
Bgf1w7W0yhKGmHSx3TxmMfyHVwjFupf10ZqaFH7kI+kpHuAiwJgVy0X77UyQENhD
jCZnO0OgcK45PkslIMOxotnE+wGz4o9UStOGkGnkLWvahPBgYRvdJKrs4B6JXb3N
b/JMiuwqkOKjm569f056gZFrVVZveWLR2yKNUM/9w4hi8fndbOJxPR14E/0BcpUL
urVIGhi0oelx505eACb5QxxEAy5CF5oWB/dlELzWduw+mVYqXNoKAr6zyJuToChf
8qmW69bM7X/0CZ4hSFX34RfpZ+cAS30xs7FqwBvbDnPXZNuFtLbOLSuF5eSRlzLA
o564abvFrbbHEgZ9nYAsCn7kbEH4RCFadROfFs8/raFk6+QYm2YjvSE4rdmMfIWg
w6oHUuen+kmgtXNBUqIP1Bm8jKSVVR6vXcz+w86hXQDRlNA8PNHaHHrRhKliIRJm
kt2Jt0EaTmUhkzSonXIURBbXVTAWjxO/hK+Yxb6C5EMHuGUTLS4upvIal+OpK/hP
VX4eF6xJpxbh/idbWkZuKKSNCJwedi4WKCIK7t2180QVexwID2SCeO1gB0sPGLRV
zZU7o4Rv6sS0d41TdesUcxRly+WXLrYJ1uctpmTEVJuwlaFAzerhBmF2YGut8S1B
LAwys0vnfLwO/JPMV0kE/ecL1TjmoCAT73d0v9krjwZj5yZ5WM6ODT1Lgd3G37dX
oSCdU4avKNklQMNpQz3eGP/h2pmR+X8rXb1wuv+KVeiQIrhIw/a/6j5oYmS5+6Qm
kdNg3Qpv52XHrbFP6WlxrxKOGPOIbr5h8E1Jy9XUnl52j08A+aRKD/MhHorfgVHR
zmqoEqkKwsDFRiZEr/ho/6VrOCOmSKFmJKNtF+bewEgJL8/DcOHg9wI0HUgVYV/t
riOBB2F86VfbkEuSYlxWu5ivmxAZHFtxk+Zqgz0QXKqyVx11Pl/IcA+HRfU9az9t
PmnQcHLVgit6QkgYa8CBxeyBRlfwo/lo+9GTm5su/yfDd1oTfQF8WiN5zlN8d9ze
OdrHIIkuOGR+FOdIEwC1/4Hl93Sf4G5QWolFvMoLRqz/r5HofRt2gPh/ocM8cMo7
KKu3NvrAapLeAGdjiIqdEoHaiZTt37rbVz3Cgi0GAsRjbf9mDYT+EmjpGLec0Yrc
e4/txpmGFW7sjOSElG7c+iM0HupsbzlbFgbGAGjqHwxlebd53DqqC7V5HD/WC6vm
+fDqv556fFczKEML+3+scYcg44+KV++fqsjd7aTwFXWi4RfXNWL5HmNvLukkavEA
Al4ECUnOexqHvu+O+0Y0rkDWViZkzBhxGhLptbvfy4ege6ytS+MBWa57Py+wK+fa
Gqv8J9IYXEzujoL1jUoz2D38CQZ6sTdlNR/p0veYz5gxx2BIYdkUy3KDPqH8/PAd
JDnYptmGL0zw3oGgz1uAJXoym/9g4v11ec1ZfxRCTAsJQ+L/mZO/VI8LWjz5cYEU
jXdV6Xo7dTOLenvv/H8evqwX6g/BK6kbJPbtX+wUzk7/JyWDi+pKpQulvvEYl3e6
a0TPLJ6RawfvOPptF17tx4OmFGZxYwGE2HRNjzZGjiakxEBOdLc5nqX8hy1Y7Eih
5lvYD49FxfWA+l9lFAGDogI6OnK84p6g9OPwA5lxJTT/FzvN+1Aa61ebPX8TrsLv
/AUpWt8asfoBtODm7HwpGONt8tYx/+qFaeExFWLoctU8i4dyxBr0BeQe0q2xT7k3
edY6UWkKcZcSu9V4s09M9NtHfC4dDN4G5ThJb/VIrhuP8kAFYNDoRnItg2NfREDl
LiQjqTIqYMyyQlrgAeHOHrE+oZnjHdqlFz+OwQ07USoRY3yaeaTCTYW8tgGFCRFM
0JmR8LBDQDzX2/CpKNkvkltD35b4B0Jn5+ID2SG00JnZ9ac79VHu5Ru/zdYZXJ6f
Znu5wTk1MoRTFZOqWb65bwoDtyq+xOmYHZrjOdE9+c8ZPCb1meLcCt7Od8khHfVr
SQQl85PwVVpAOVNr7hsDBYnXE4WYXmpvtL+eBbQMKAjMa506mQPiGtEZhP+BT7h6
7H58OgJdHpbQYwbHRgbe+ME+I9hVpEHqjHOspwr37Dy+yWYibsith4hbM14Xkuhg
Kilyy+cBY3mC8RHvBJmYPjFa25McmjtovOGhtyOZXjeEbTU6QlaDfSgBBtLvna/0
zeP99HTeQRveRf/Ro++kBAs8vV4fdlWiRhVZWDxAHZrtUX+fYKXIHtWoO+7bxYC/
hAkE2kd+Yijcdgy+aoiulxoirG3Ilo5eHB577jXNdNtfpc9Ejxrrlhc2ekutWFRB
dEJsxLjnXX3/PqYDu9oIHotqjZoc3JZVidK8mPUg5afG5LhPDS02usg4NB4q4Ec+
asSdu9DBHdWTPJnyNWvkjdwbV1w+MY5argDH+4sb+qVISVAS3+ES78bCqxxRJEZj
aWi2L8G5AHLbFiIV28YBKCUwZxhGFp57EOE3XSEIXdxIXDXeReBoQkxcAqYWeMv3
y1wI3mfzZ6f5VwZH1fGCwMF/FzklihPI22uN/f3OI9qqvOoT8yMHKD4QUF9Y9el4
N94Z1uZkkOiyxjMzIsXdWt4K8+4iLYABN3o3Qmxc5HJJuR1z6lOFCwflXaNLR2uH
YetDq/CHSB3LrghDI+xU6h5PuVMXPh4wYSnGXGSXuhjXrLNBv80+dHpGMNeDU4FN
+iB83Ko3/RcScjVHOAH3aw3X7FYhZdJEeLg2n/zTdssmHRhsYHa/D15gPz0oERow
oduJpEyhmcAr536mbRSiJ8Uq/6uxbvnQzHn0/uIG6E8frzryiTNopwWDt+UOMhrL
veAXcaEY36+mC95HpetRK8A4grfwPmPe5962jkP32A6yEWvWtE/Nxb//LxgB5bVg
gbs1NZQ5vdracAevyTBQgMPhh6dqXZDfAIDafGW+GB4nhv4TyBeNS9PB00tMmSql
C9zX8/Hef0WY7nXQ+iC4GaTWpeNrAg0QrbzGP2losvdSxT1DJcTU/uqd3OTYA+xj
DfZf7O0hiA6uwVQqJXbmUFOBwenOCGRrTsz37bTWUTuPt60HiQF/xez54AB7+xgN
PrY6/AjRqI+k+E5rJSOWWLJWj9v9BltXwj+QnzgDmOMuA+F2vQjNQIrkPFv83BN2
1Fsz0DCgcDsD5emkNNBZ0NFz1sd0LvyvZUaTygx7IqPxCh01YkcjLQMRZT/wmo9F
ocP232Cbmn1WLoLNME3gMveow/y8N9CxOz9AeCHZwISIhZ8qJ+QupKprF9ROezis
SXdrPH9nUlAwSydHnsGRSy1KfhjJJcjv5Mpkn9o3pl4EAPYTJpVgCmjKwvdONmBz
jYG4E4Rk5IooAWRiWsjVlVYwx5w5Uj9RAHlj6l2UFX5L8v3qabxCFxHkIHuGO7Dg
FmiPgfxnAMrfmZ/QquoJoStqrdENscU3wJeriVoUlZeglAq1wIEF8OEn3UlUN+q6
jyK50Sg3+wpoB80mYWx2fTYdRk+ql8ojecewl5Zqhh2glORemJ1dsiO+QMcUn9+1
7rWcXYaroqy1z5eWEXKiNAMT21SguXVS0+iE041nJ+Wnvwu/YRQkGc9ZiJEI4vMJ
FWCom0TH3BhTY/63GubI0UU51Vz7kVxoET1W9TNAE7bJa+W7Cl4QvuYgQXJ57hnB
4prTiTNi2e5PcF/GxY4CT2nRdzTNej0WRomf/G7XeX7bRHPdk6hsJ9QcW98dOVUw
+tFFa1PA5PTL69eea4r5K6bSeC3NHZAzqsr+2cW2bKug6Fee2X/G9nUBF+sSCbed
pJ9mCwrdjS+j6sswG0pdkJTTaJjJINRPg9IIRA7/QoOa3OOBhCqbCvu5sGttU05R
n8zQ2BA2nr6frYD2S6/rab5nnk4DsNFKKUi6KoCJooM4+vOAJo2JoQdlOjOurgjc
OdsUqV5NCK9XcHSL9koQNQu1AeYMd9klLaLDdFLMXRRX2GY3DCpjrwlrHpGPtOmE
SHbzp8dO5BRpkUJRKinX/NnB8pkEbhQiBl7AWlJkUEYoY5ZuSljlo1RKwE6p1a0Y
MZY+Jxxyx8Ml6EA7Ki6iC9fnviaMKeuePbiJ36GuuRmCBsXpm/WADp+8vPXN4g+F
KAUC+koUBQw0PGMZkLs6f35SKt3fJsQEpE0OE7U0CKAmiAvKFlWeYNPHF9UM8UPZ
mDfaoXoIgFjLZyfoVfB4Ziv5+A4KTslHWtbUtNJHIvG9zMli420xjoQDlpvvn6DD
FTSuN3yd1/ohHjqYiiXyt/RxGwpvxNgIc07HLlzdgMWaegk0JLTcKJz38Uz5TUfK
5pCqZKoU57xZjdV5Lq96nb/KHeMEVDUy7qji6aBv0yu3S23S7iXl4TUX/847/5yM
0KChd1zgt7NM6QkmqVEMmskMZy9oI+YQrMa2SjkWiLGH2g9kg7iRqtC0+LP3QFCv
hqwGMNYFJWPXFv0/+4IW7mCA5CshLeysvWTjZziuAq1JL5q1ygf8u2zWoUeJ0f84
p9tNA07DePgufEfYCmbzgkwo9w3BDGFFVZSS/NG9s1rgMpFpsoG6lnGboD0R/QrZ
qi9MZxcoZom+GYzziE8n3knG9cjRrVhQGS2tRI658lMVjUh+0krTtbpKixfOG97o
9FxHhPCITD9N1+hBxFNWaAAzTozk0atVgX74eT412Wy1aIPP46X2wr2QRrwGZP+C
ysWj0DxKVgQbeFhlXgk1Nk4DqolAPUAdeasLZg0KC9/LjUTsAZT+2Qk+AtIeL5he
jsPgxdgzi3Rr1cvYkxEsPfzg5lBTEPkHsEGwmSsQOXx7GA674Ojlm5vMSgN8t6WS
VAFlbA17WxzochIJxFEAahpZIdtBiyjBhJgoFm43lt8Q9ZR0nI35F60pIgBxYGyw
YxLhRsytF642XEMiucxzTfkdW1MS6SIwUkR7UyndZHfIWsp3CH0MhPthSjkUE7Kj
JOaBA0QKbMfHOh/Uj2aIoUsYGWUepniBYVC4WfFaCECxWP5v/iR1wwdFyk20s5ai
044Do4GfnmWsSg1W7dMQ2Fgl4pOqnJHaCQPnCZ+/qj6Hh2nzl+zTiEqJNP7Bh3Vd
K8IY7OqX5Q1AyRiEEgi5aAUf8LXQ6f0UvFvR1++n+wTSk0N6znUTmz/U9v7hHloX
o/qaAwjkNJ2dt6gUJwVND55lmwMmHl+0cNM9PeoMJLenTpAbApNV6QJSqNRRzxJ0
DhGswT4GcxQxpH4WDExaHY5ZAlPPWoBH1J0dS33YZzPw5gn13IY8UXUzDR1sstTE
nDm+lds7snoHrqA8qhlRN/zwdvJ0tELEFHV/zlvls/w/B3kHWrTJ1eoMqCyERrOY
gMiAFgEYTkqkbg1GeTqQDnqFqlAsBO4auhRfYm5B3IJVMA51hnnDzByYtcg+N1U4
WzBPzjU5ZPv86K9xOVzX7F1CJyPNqLtD8qoLxxOk40Qs8MHf7PFpIaV6f5iP8StU
GSNIpUAiMew339S6NuONsIZ+Y3q4dg+Edc4hwfKYj5+JvWLGf7gDj/9W7zhtgzF+
kG3IZO+qTjXbYjOOY7BBqwQiHUoaLs64bnRLlfTLFbLvf0Q7JShJpsiY/mO3M1LA
muuudme4/7kxRla7xk7raGx2Lt4XMCleJCFt0lQiCTa0Riza6pxLOBAM5y9Zo++1
ftHFI9nYUeXo0qrEYUdSEOACLyV2jdAXZ8CDHa9I6aIMLD3GjiQP8/hH3NQCaUuD
3kLfg1aVq6PbjVJCt99uuG9eKN1QgDVkwzeugwrokq85FnbQmWiI7en/bx+iRWiK
bkOjBAaf/nArmcfoKf+DsvSULN5pbUd+c12yFnUEBGJfZ9rmL2RA+JI7K9Zuxmjf
g/7jyhtYNrPna/HQ9BTZqid4qB20N0yrSpZ2aahgc2rLs1Yuu+v0osVahcQ5iZ9k
EqSbbL9dN5rTuntvsideMGRrM2FomcNotfNYGTl9mikD82Sa/6Y8J4PTMQERIBiS
1B0DQFozITvUZX/aMH9Hlb2ih0rhi10uWWg74jdekqCEyusc5hdzL+dISsaUMdDW
etprtq39dFqHcOq76rpgYlJ0HsqKD3nc6AAQucmpDt9bDMHiIIHIkmGURcNQJcd9
6DlRNQerDga381bEESLUGi7QsVzz6P9ufj2kBkHaaR9nrOwY9Vp9taM0OVuQZdLL
CDhXwx19jKvGMjkl5tt/lh9n5UJCqfQop1MpjVA+MAQ6tiLlvr7ntLy001TdJpFx
cBVquXnkWxfqjtbmifBIzJCfUsL92S/Tcb3B2t4LgtpI13dKjsSGZ2bR8L3nmn/P
8OVrihfdoDZ+hrpUXoRkuYiC94xicnuxguTa00uzytDALZEQ2shc1mgC7fj4bkOs
R7acV/1AMF6t4mxGIYb2sTFgQ3bVY1cjnsiNCoVWf+k0suIH/ENqdwDO3XkeretD
IBZJa6PiiYB3qAJfeC/20jnX0/TV5qJpXfUmco2zt/pj/8vZb938iTBVn60eQaib
bYveWSQPc1c1mveJNEsjxNwgxrKzOzpC4nt+08rQZT1QZUiXW5se0stm/UA5e7Tj
wvlyLyy8jwHSVBfbPKqt8fpUrNDF7i7DVWjgKWC+6C8QQEF8jrrMxara9XDhhDGG
2PPco9Yhq8Ru489NjsGvy4edavDY0yU8Rp/AJGZgIT7koqFNXQIZJxIqGNO29EdH
oTnx/7IZUJ0J5b6jR+3ZYtH2VCUi1ZpLK0hOMyPmjBo4YoVJZVJ2nvqtvaA6QhHi
3dP37iXbHp3WWaLoDwoTwHPQrWXrj8DZIv2YlUt/3T3QlMs/inFdTw6yPV5ZRM7c
yLXKNi/M2gc/VdiNY9E5uY5kW3WHR0S/BcXkkPfoaUDXH/wLl+ValyH5nmwaRnRe
IVnOcQAko/6eCSSdY/FiThbVwcYUmYxraZunPyVHuDbVD3DVky6POu0/jMczXAk4
FqdakLgEgzGpbBgu0rkH++Oa4vkutvJxfTPdJD8j1hZelX02GEcJx2J69NUi12NU
6xKI7glIUck/LpMKMiqQJgs1cGuhJNE/Ir6Oieg0rapyFo/d0hGyz52E+uy5PA8y
2jv5fHg0gERKvlrV+T5Ajr6wS37v/PmGGRT3GgTtegj5pQoT8pDl48TOFFUHHrY6
WJKtds8a6EtuhN3e0b6WmmpDZYzl72ZMdqr06LkAH8noqw9ltmdjNR1DWaNpDhsz
5ey5aUvI6Rs/lFyGV2ZD/B5d2BQ9+VlhLUhvt2fG7sbU4+pOzXdEuNr+aJ8+AWsZ
rqrZoC5dYsVBM6xh1Uf7/jf8p7PaAaIRoEwAIfQLEp83SpoATot7fNA+H7YfD9iE
YpnzK3gRo67FfRnISpU6ra4d1GG6gXmJPsIyTrIhD404knwsStM8/By9D2nlbg07
eclRUGNi/n8OwEnt1xwUUqZRkZtOU+HmitJPk8tHsDoAK/LhyOxa+u6c9cf3vKcH
8/COrjfCADDp+EEVJgkdzbowqmtCxyhMi3Q876fx43lX8ASKZ8Ap9UPLJRL9oSp3
BoCvNJFZtY9MuCUne6D/E+Y6p+ilAeI9Oo/E8AeSDykCCAjwgDgHAadyS/hj/yUt
ZS0fTzLZZDNf+/YRMkWPlROlkJGc2WzvDmjivrHgK9NmLi5r/Ux11NETIIXHIg9E
Z+kr66ppAMtHEcmSOBVHqIqyfgwN2srLXy2cNp2e2olsp6aFHcaB5iKfPnJ97Ld6
cMjNirclVbpsAoMd2iIYDlRvrTqYgdeK7DQoreKJDt8l3WWAqYOgaeY1Zz3Ujsrf
0u9o8BI3nGz1CwDgzv5hBwvO6fsAVaINK52jMFcaGMYztctizOTx33kPhIUmgZKl
kHuGnjv4AOHOffJFXd6XXCvHEvPg9L0Kh4Gs+kjUXQFvhLCiDv6qIuhy1LoY31Gg
03mLGrEwVdAspOpn+W0LEpFNtkzFFJCVQ2sgur+Nt9tJxYJPuaWdZqi6jCyk8QWg
gNGDkya+FHCfqZQWksEy3KSxWNrHTiAmBvWwSGFa2l7usuwuKdKGCR0hKyy+mH4Q
ccKq0kw0YyB+OZeE0bPSSoTBKuUCwAYFTrx+UaYmAbnVtKyzGeXfjsvp4Fetl/n8
NJJmZae1Ig0pnoYXqatmA/+wOjmz+LTGUwwrC5MLZlfDlUPlkBzRF43hcqNW7bnS
FzANRtREB7Y2Z0Hwb27cYdMhanzv9aswKZflbXcEaOPBWRWiFevmnq7cW6939B15
8m6bzqGhtsZPj0ELZ4vNsxA0ORgqxDmYXy+9GaVkBgyEbyGL371sDhEyhcXX7iVi
aAdYFxKWxLiLt1WyomwXKF8KIa6IekWpTlWPUPqB+xi1du68Ss146HvCSZloNnaE
tJzFeqJcJkjR1NeNLkkOD9jHZ/FvnZXrtU3z7qVrtn3Not9VfXJv77pRx1iISzmH
FDqQaUNRHR1qFnyplDI5DX7IM+fKQO/8OQWqvWkydUhkQvBHszsr0KM/3eK7qaFL
zPIz6rWkinNZOrc7AZRzUY/aY6zk6liqiLhlUbx30SYpiQJ3xF8HX9g9uc9zKmD7
QdJABfymoReEwGnUtHph8dSVwZkD9JRdJ+3X0m1AxRwqwDCKv0+0hUFvBcTzs75E
LZvLBqpFd2958okXpelqFMKB2w2Bn8UB7h6S06hhcAa7zKuu/IKH3BhlXPpj5Fpq
cLlZXGs6Tc6d/gp7DSiCn5aHXvuOlwm4i9upSEoOPBSd8jHAiFnCj8ZQb2A0Xgzg
hLYbFdbnJBwRS9N1wJywq7BO5UhVn5jUvarKjpJ0Vx4B0IdVUiNJ0kO8G1q6E+Gp
lIPTp3+yF6WQ2FxtmyfSWzd+yKUq1iNIV8CWLNg9EPyzudjgpaT9ZZ3mytX+B0p4
XLc58qKLiMpmmT+9M5/wxcFb8m/guoQyuowP3jwWGcmqI1jL2Lyecj7RQTNE1j1b
Y6nvzXqn/cddV9hUlihJ43SG3U0W+w4P/gnY2i7BFTsYd3DO3jqUIkOtHmu2oBNv
Pr/Y2EfoPrgWzkMVMAZ77t/NytRCKldVtMChUabTLafTX15vcoRm3b2cui8bchq1
Pltyktr+M9FdNSr0Us5y5JP1YnskFXEFyoB1S/sodpZCRDbYHJ7s1DNKod0cZbYL
HMVQuTn5VDIRQsyPUwDvkZl5UnmbHHdcjP6ZnanwASzEgGDRqr7aNj9TlyjpzbKv
1PdowEF1YUGzOxhF3+PA5gjR4cbOAnfnl2rvRbqy9ZB7zKhgmgoHB1c7XH7JSJlP
yzCHYF7sjqa+kh+S1hzwttie4lyNOaIfLNEy1dZec4bfcNZcjVqbsBnUyXMYytS6
8moS2D9NNo9h0+dtyZqxqJOUYY6r8UTJAzSsJKg4mMXcUJg7j6qoG7Vckl4WJd8Z
IydCPTggGwdQOdkgTfZASkCCv4x515M0sERxCvsXWzaycSEXvGT/OvS39yfn6sSZ
4HyP9+RK6y+don0jIauiu1TYecIXy55pNSiqAuUOp0Ed2Ht1JUSN1cpR2WNg8UIH
5XxZlQFlVDEmZONcN10n+rTkJ2K0P4CLwUJmTTmL4JkgV0TENo+axmkUoEZJcLZA
aszxyLHF/rFL2DE4J+B5YcbuxGw80A0ibugjJCb5wRT6eeQHxbTEZOphCK+zYUxP
lUBmFBAXNwZF0/kErApzpWKnYdY9XcwlEBWQtxhQayTY0rTkaZdmibr3LtWiD06J
jM5PI+CnN3le2SxRJl/usMkzs8RtlsWAQCwYytK5BKZc9RJ1cXKvgB1Pxi/VU04B
XSBDaUGd1bRXUHokOsZPl6RfEjGrGTRsVpe0AOb9q1kJbmuTcxBgzfARy3geWno4
sNkYzJBjQ7ItEc+YNF8a5+4sf7AOpJsJLgc1RNQc6c7r+xqEjejr89Pw7KFzoPad
o9M47wxg8z7yS0A/pSl4Fe4SkqtW4z3aO1Qk2uFShnuantdOOngsdOHGxT4o/xlS
Z20PfuIFztUJMSNqFr/Pe+wSpVn6Cj7O/2P7Wqii5PH3AehOYRNgSNpVE7kEf3u8
iILu6HBR37YwwNZ9IUILQUbLShEfJ3h0Nz/UqbJYvTQ7Y3o1GokInHOMxBNKjAyV
+laM0b29fa8poIybasZJrC61ZIF4UakT9dq/oehoYd6y6xGlJyYJi3zebTm9N7in
flLsNccFK8a8G6oScCWJB1U7h51yXExpjMK53Yad1EgvcKjZcLs9pr/LCKf4qvIy
dNFxWNoe1y2CJROIPxNe8WGTUp8k77uxcSgowkY2FAZinSVahcaKL7V+jYRupKxZ
HDEr7bUv5gbv3aC8y5yKoJRfFbVwNY3oWPPXBBn3U0+IQA2bJFfPNY0xaQ4bTOYr
tlbNPrAtIjKXy9jnfnBWtOkoHr1texVjp+nod7CpH7CXRXMEq8OgWTSfw+wGAKzf
bSafz6pi4WLIYF59fJymMfCC3JddwLoLWC3RdCZtuKBx9lvx83UnxaA6Ba7KCo3B
2Hau9+CPyM66BUMykS88T4lBNIAFF9QG++3RDt5YDXJuOp6Jh05Vaj6M+AN+2pmQ
fLi+AbYkpjASuZReGv24qmX01PMsyi/9Yd673wWbxkpwbeYUvlEzwP6RAIUCd6Jl
FiBj90h8Osw7utouEsYFHlpXi7950j8vZhEfmfOqzhKtskZGJlehTvIObymMt+b3
GppmpPqftLEuUgpjrbRkVukAfzp+z0xRelvB0W+VKXpAwX+4a1LwZiBt0ofDQQer
zK1slLwNfHMfIhD/BvTsILcAOcTgNQswXb3xg+V9T7uIpnqZxo5CEUpW7Ei9QHtX
qMVaAtw8FYbceUw88tiCPjJ0qE5FVXWzrlEXthAl2+sH6Rm6AKXKpYOKrUPQ41D0
E45fFQhFhqq2EeXwDbCSw2zP49HLRGvcOXbnj4B9CHqGDJMOfL6eTCJ5bN6UB6pr
zufx7jqR+wO/634eJs+OxDNEzMxtOFoaCbB/3R/DU+6c8OY70hiSm3fb+8wMuE+V
adhzP1YhHsikS7MAk3OAxUjnI6A8kxd1uzngVjN317GO9WRy0BUrPniZTLY5Inx8
ZgWEiBlQIb6UtzgthHBnrYzlx6uCjnkA6akxUxJE+8WZbh0t70w3Ga8xXLA3RkEn
fGd/HctlYdseSoh0NS/JsfvDKzRTQOWFp9PNnIhat3KoFU/APktLtlSDRwCaAZNv
gWecHKaDT25B9U0XNR/X5KHFeKqA6VF9KFx+DQ+iZQLu+f98wJ8y8kto7lgrHj5j
h62IPnTohDUjiuvSmWRUys8hDZO+mF6Auk+RXmA9q+KuUFIImhbpNjwiQNwhfkYB
Ak5qtfZT2PM7442SN/WnJvfNhDtlYNgfIhRsKb1phdED5Nkjif82Cawb1/6pRYnp
evh71YasYNPEnQoE5thyLZjSlojHPNxihi4QfqvJvEOcs3stuO3jIqWdfkfGUpJU
kikuSRzI8OU2cG5KdP8iOVpckS9HnwKGfhdjuXilmTizNLm2Lzl8/K9ZhKPvPKoT
yYCXKmEuCoNFmaDpyXDerDEU+JGwjJgJffYm6P1QDYKoI6JQwh0ks+bxBVA/2qMR
0T/InRFV7cEo7jfqT3KgDyY7dNCRado4QLPKUakhRBNi6pe5DsoCtXQN7YYi8dVO
8bHFM330E6NQupIOkD2ro9phRG2dgR8+DCmbYsz2OcxsPAqtez0mPSFdfxf7aIOd
A1/Ycx/wFjdXjjnNv45luXBwwXU9zsoygdpEOe2Kxx0ayR3pD3Hvj7sus8AZFAo+
1d0QOCuJNYkoS3oXgtga7/M6uWX+yoltA6xkIH0LWs2lcYIoUxOGN+BmfHUieiPo
Pnbhe25AXUmeGu7peK7gS0+bkHFScFS+TlqWfZ0IN/G0JbCCyAtRyloE7r87PrbW
dWOmSrdmmWsEoOskj9glDFxIsWKt8Y91a3cbgMIz4kgXPuP0NoYwgpL+07lyKh07
dK5br8EyZceO5k67IpUlJKoxMREtX8QLktiqjUwOoZYJvN6TIJtJHGZwFjNmYrrb
TryUhYmR3n9yeOjEtY6qMHlPUV5zb16GECf2l3in0Mm3Lv764v8XDtbnjRPKZe7Q
P1rZnCD6AJ327Z0KTcFTskq9DZfTrNmGZHozCSLaXelCbWJSngWwz/rGRIuPYNOm
zyfREzhPHFAQm5KoJ4b9PQBFbMBQS0sHA2rp7GwakCCKeALxid0LIJ9ddAu8Nx18
QIQlPxTOnojGeMxaRCBFWqOzcRxnT1+RCU7bCBBgB2ApoT3oXIbbuXJ69aqgJUoC
KzTiA30B9oXV1vXlcYDG4frRLVhlDDpnpAplXeEg5NUwLwl/KjV4DVfOMhbAXrSA
GRzUGCiidSNqdDZI5Y/6gRLTDEfJM5NLhh77uLRK3CnzEotxT1b+MW6xmWlVSkSX
5vJzBFWsSiGYkxSoKJGVFOnhkb9mLt8yWKqH/9plfX9BD9xzyQRqc/UduYUYa+tu
cKGabvje0YiImqJutKlUScLGKA4/9/TIBUTImXzh7ZXpD//pP+hM4SM1+VUcNLMT
eLcBkWHxhN+kYJcyGjrmDS0Pgtrvb238jHTnuG4KsxLlxRWpuO+RLnbL414ySyjU
t0yNZX3HYZK2wBkG/Ja+wcaVMKXc4JkTPlt/9EQek1fJbOdyt4PxUY3BXgRlSm1r
H8kta4jIFNbCnAY1jDHR/XXsR8BxriYYScskHpG6mJ+m69lAWjz3PCAkHvvOLoPD
PKYfXwDAmH8qQTlavr4vqg6zxRPOGAngs5NZ/75tqe3Fjmg4O7yL6tOxCy68ikRz
NlD8bm7H1rpL6axn5wlkFZQdA6ATvntCokFRJxRvvNG9OeKIbE2CqLULVKeu6sSe
HDNy6t8afW70CfXdFx1U/it1np3+EPFHJQUbSmQp3LKVEPjojW+RGEbCFcNIe9kX
uEz0vMx+2rB00gv+rbYtBE2M1j3F8soGMKWE8jt3IJoPKOmkVxw0gemOepN8o7/3
4Bsy2j2s7UulYO7DpfdNHf7M4IxbOnu41AxqxVfhVgKlkpg2DLpvqfUplzepimhm
JLDbcdftvO954xY6GsWYq1FVjbu9cok7bV7iFMRFnLrwOyGmcANYuiSTaiarm8Rs
DV4nBtciKvTy056gI4Kb8jvljP35+CF0min6950RylO4voayInO5Wqcs61cS7Dft
6TUGMTqRTi548F8woXeinKbBEqKCah7FL7mgfpVWZxVeNidasGW5o17cjNH47qtX
BCD3I5gjL2C2xD+LGuHK2pSYSD76QWm26p8VkA/zqxRSv9YNV6uEhTWM6VCrWUP4
9Tfg5bMD3WHh/T/KOfeMF3BUnJ69lrnhZKWqm41HUT7pBSAYbTLgttSDYYHkjA1p
uCACSyYw9TiQhkHGOZ2pVWiHyuBM8EN/XtW/NX0Y9sVSWVcQiIVEIuRNoXa4xYAy
fqO2CnPy0aCEGfy0G6PBfYb+AoTBLJKk3Sv0/mU10lNZ9DKb+v6j6WtVg6QC4srL
DK88FKTL49PMF4gNMv7gLvSEHI6OmPXXXeoda2L8rwZClJV5T/LyN9FfYvL6TON4
VOzpygWVnjTx3EaIgTatXsbUdsqR+IKvW0py+8GkJiXg5rjqNULP91mk9rKXTjLm
hVT8xq012+vXOwEpnF9HnIbNz5QBzLTk/LOi9gg2TsL50VD6i4znK1DlvkjhTOKV
VeRY5HbO6+kQuR1vRnc5w4Mc3jt0UfOEaNMcoZonVQboaOBp3WFtt8txLXoaQm4u
98vSLgQjaCzft0yDR9sRth3kmUT37Sh7l2TebG5+Up/CDOWDytqaKndIioJG2sNo
gyyhf+DdOHITpwHYFEhHw+lCgpiSgvPpmR6oEyCUagQ8Nbf11dLaDqjL77EUBqtA
/C3lsCG1V4htIngfT/YrQ0AgRzxt7GgKUy5okSdSsmUhTmPMjHdjr4P4UsicFc4m
5hK9f0hOwqyBe1NkAElfZSivVZz0xdICCqGM2YeTo/MCswiPD0TB01l7sJW1+njV
zv5yhWIsq8JNmgebUhaElG4U7bpg8l2/CBnzrQmYeJr6q27JANjvGcBmo3z0FKHr
jRIe4h70GD/bGmFMK9c4LsgNko5AEnCb5zlte5OPTYKEltMCp+ko85VsTAvj6iu+
87owKhi9WMWRiD5lJ8p4M3YPazRdOuSBhE8rFHW+anAkrfNpR+kCdulYjtyumYNx
O2yWkatE5+/Q0WkO7Wam97CRgRrgKCUj0tCcCd6GiCWtRP8JMK4d5NA/UpoVML1e
3puoSxE2NzprTRNYYK7DoBNPechK/MuMxaZ67EKpSi+QxDsFJDdYl3WU2tAHIcU7
MQ/JS134hp7KNN0MyoA2cR42JvKi69Rfl+ErdB67h2bNsLrWsyBVuijqNiHtEnNS
iOCcI8bh2JK53yBfXB1RtANxlIxoN+TPhbbQlWp9gGfyV0sHdsr2/87iP5TppZwb
Q/fRwthmGxI89V4eLpTHTBMgKs7YBH8VOsB8DQ/lYE10c6oERmrOIHVwHRZ1Llib
4DcwuJHcS6i/lqquy2x/VmVAEXDKsm1J2YfabiM/URn0ec2vt3969fBq2ItC+XZZ
uqHVacxeOvs/giS7Eq2eIJXC2hxTdGur4a0MJH830Xc1ddFZXsSbfaVm9/DxTk3y
9CqWrbCjM21oAOSVMwTqUksjIr1k1T+l3ABrC2m6G8pvu5HKKvfTfkIhAaYFMAEN
OAdq4fEjOZb+XWvvIM19cJivHsFYW1iwaQzw1KGPGmOcUxuf3OJ8tur5NTLicVvH
6KBht2oSbfUbYIyRu8f5hhRkIab3u18fqEWxo5NHUlPLg8jrUhI1S8tOi3RIxVzO
FNrOGOsinX17vb0XgXzZUNGdLjQZ4TEgJ1embzgWpp62lS9xZev6QP8W/5H5hejM
13arZB+3SzNurdAVesDe7GbK3RB3He5ssWwKs8FdHz6Vre3RaJL39B60rF+WF983
ec60BHF7dUsTazUgsKv/dfiYGJ8afczullMa+ZannJYfHarwcPsU7NR+mfDbDLj4
cTR4oxVaB53rAM6lYiAEXz/nuTzWbB/2mL9kyckDxIigpOtQCJxczQi2eD1ZtKZS
xMN0XusOi4yOrpWI33T5uspxWr/IugHBWwOqle0I9+i9aXA0XdUPySoG6T5SGOya
YdFxxOIZm1U1dcJjrVT4DPUrlsOOW2Ak4k2NtjsSExMs73bGAMZzI0KkxMt7fPFg
TwFVf9O4otaHvoHnJGRnE/RWnGRlkKcv1+omUftWoBPo2BsRPjj7ljjPpweGJ7S4
s5V4YzTiMvO7y9b/A0h1+7JWO4E+Y/18F2/hAWbl4zeyFv2SIr/LXYg74YD0djmx
ARE6VoCtg04j8dB6520i/dEBAe/Feub9okizx52ZeiDPV/gmOl/+rR5PfxOvk84C
0pd9z9yHAysH0AMeUzjHITLPzeC9H1Luia8x+qCPtap2nZAM16boMtT6/yCFIzwM
ixXGNzqVDKqkX2U4uPxeZEhmfPJR1vokFI2h5pfnQ3NGxmmxMg+WUGTETm9nkXnH
soX5cVzuyyNF3Qdt0VUIRlZo8GIn8/KYLtvonGXz7odQS/WeByB584fnGtZ9GzFE
NsJn2QBjJuN4Lgloj0K25M1bs6wBGtfYadzajcKWrhUIQMqNP4yGrJUcrrGTJWKy
425eiqiFEvDool2KSh9DZZZylZ/LSd42WCvok0AqLP9vP41OhepSS3FS04kIalSw
Q6QwclQ+jeq8EIBjf+Alsh8m4s96XJb5s+7RxI94qQgAkP4CHf8ipJ4x4LJxkIil
ZaA8TWPL8jaeQ3ofC/CTqGkNZYZTfqweMpNwc9AnesM9ZEMS/Be5uUDtLWHc6OMy
qJ4OBaEPMyzAuHnYnagcRXR/qALnmvKRiF3C1gS8css+2/ka/NdoIobC+QArKUXP
00CCQhgYZxRN5Kg9Dz/21pBl5+mpfH4cNV6JgFqqNPh8XyKGTdGHQ4h+wODLJQLX
Te5Ihy59r5WpARk4a1XvQSF5fx076HX/mGk+47nncw7OSDLWaNX4QJZvoTPusIMf
Kk6qADtiMFNy6MAbUEvEhv7oTuOrqn9LFMiQF4B5O2KBWcVN5x5rD2CR0DfNtxte
ruR5xQg/Nz0XAxoKIgH7e7SS9ektUq+L0UFb2l0NBL/6EYia7aYfybS+YVaXBxLr
nDAr+sPxUUvQuXJQWvJYkpXp4ASyv9o7ign5Kd22QnJKJdyq3IlEt1aD5BbS6RmP
L7kHE/nRaZQQpIuba6l9whthn4ystn/GjlzUvlUYui36KztNpCrGsMzqpkOlw25h
otkeBLfTB2t4/13u0CtgQhtqW1a8NhgIk+cqoIy8UJvaNatpJ41WvWB6Zg/7x9b6
ET0gcNKEOol5jjFnjsyR686Y2VzlDlUwA7BH0jnYjHagLwJxzg23hEODdBFBykxJ
ons1kt/tqGrsYxG2pHaNND1Rmz6o6YPx/T83GY0WzWYqkd92HJl/fH/uV3Jaymz6
PORh55u7H/5k+rL+NelWIOlF+KuXhm12mJx+OZa2mfIFguC4/6GYDdfVRtR5hhX8
3NcGOURk3GxkhL+osTWEMcqwBd1lBZn2di8M7DtLXD8rpuXPYzHfMfZIuqV1bMk0
oCOaiHpP/8TAKb4FITSrYvad/17ES6g4DV+9dq5KHG7MtTlDRz/JKl19R7QoMiY/
NUAq/m+X0JC1qBIlY3OVTZg9JdDD47xQhzKlLpR8faum2ZXIt2lgYMCPfK9FyJZF
iCiAM9vtdfYhIDvUcvMCkpVLx8U/eV+JBVHQNH8FIh4/Vgn958BLf6pguXNkf0QM
F8y2Ou56s1OYdiEfYntT76VWtpbO+agq1BwMTMPhasmJWJ4q8KCNti48ayEuB2CK
wlYnxwzWs9vID4xKdoTj1U0NCH4ETwE0dUnDQNdbNnMGX6vMoMiYmI+T/+DydYeT
eD/MCDrsNe9aGdtWNirQqDNdtOGrn5OG0n2ZQekfwyvsFjq803LfkFeGQA1qaDix
Plwce1X3p1eMyfsuMpW4MprJrJCKfZXgHmeE6brrMYeCxzXfj/zsFISRESDn/bs4
E5soYWqQQF/JQhWEUTPMmBqdy0RGJgNMLtCfAqpPmabNTMcGETNI1o2iJjq+Jv8s
zGUJVy1MgjqaMiY15fBCCvR2E+yb4OFJlYRPhQniPmqYZ/cpoXP86ygO7jAEPQv4
z2ZAUf+uOOwjJD6I0c1w42HLth7SakSkw0BsoRkj9oB98WNcmENPSSnCSvpY0+8O
PL3dYfTepYREk/D7TyjtQsQiUOS3C9VbIbPeTAOsDiFeTx5C/THPozufGiNZYzXJ
fBgMdlWjYaAI/2AIs5C2x30Y+sbV28SVcW7NGp8kUYsnWZtWucAzOMtfAzEsReyN
Kc+O1xJGjO98jHCdVyp6niIg9lcVCPx9vyqKC4wjDMeZ33rxihHMbP6A5xNwFk7y
ltsc85myGHMYrslGEDRLBc8Aphq2x6+IS4efFyqe/uYcwV5ch6TFwuSURQVsoPY/
3yy0gUCMVshoI4PDedAsuvwZh9HrHyLITrZGIJ207quzGjf56U0zyWH7CeFsJsod
06nM7BzYL0heDmZFM2NQ8ga8CBTHWehC8nwWGSHTv8gIzvw/qaLGP3gT7esLWoyy
WYTSE5yIQbljxylKaXCe2YLCPyjAxCXftgxZk4zWIF4i1Q3LJ5KnKaqoLeXBGhQT
YouyXNZZsYnyv+6lVOALnYUH4fRHEzO4Bux7E97+LbKCrt9WsfLM/ltW37Vz+r8C
C0kVPHHOlEk0O3JxlFtVnmeoKZfT1B7+WEEwrOrpjSRYdkS0u3uS0PNKo1kDlIlE
PrkMK0PAWFchrztFWVm6EUMHAfDSfStQpesp56KVU5alVF33U7x4cMv+CAJ3BC6K
aJj5Miuebj5y9G4hGohkZTeMAfba5DCyu//7OWlPZNnIV8zknAaPTCaAMcdbwchJ
TZxSBoH0tqFb4ukNqz0yfroqRd5JuGUKUCyyXfRrNuKqKl1RXNN/vzFBWIMABQwn
Aq2Yu4QIpBngGxGUnbWnxn53NMuseYpFsJBcUGHb5OxwMM80xsqisjZ/CtaPm9wQ
AKeda6APjAbG6i/YVP/3PiMJU/NLscwsqNYWic/H9s7J7fgAdo84lGge4sDACxb2
PmwYNKecbztlB6ciVFDnKHsR4Hh6oIB8e2KUJGa+YO4ZM/y95I2CeU294IY3WXTB
CztavlM+h2kSO20QjSG5beiJjmgDEvdKddw4d5yuq9XoYi9gxsX5n6UcG9A/+yMB
xVnSv9fNBNr/S1BXUXCvAhmccQtIU8rbtntb2PSYU9ejA8gJ8jUawJSCrHDrs+Ek
GOnmhtitq2N/elwtX7jyHvXoFcMg+jfqoDSMl48U3Q9FhB1WXwAPYAHI3vKfnL1d
9T9S/4lEVrBYlgi/W2cbf3wVv6CMWunb82Y4AlnCwh0+b5RQWW9311On0HVpOID9
M3RFM+Sz+SsmVNT3d1JHSL0x68uwF8ETctXSFjxaQewVf4blI1vCkXHrG3ck0tZu
rgXNA+9AJ1D4KNlyjz8VBx/3pqm9hvgj3ig0C8v1T76/plROF3Wdtx06+1BO0GAN
G9ZezLfB8Cpyr5kXaKh2tyXtrlq/xWvjzP+9BkgNZveo+G/NYW797N71OOVZcmOs
QdzF5rnWYCElo7HRTGel6KfgVab8e9I6trHs9eIAR524u4f2PKTM6rMIMttKXY2u
m01qgZkznR0/ZiaN9AnkKTOgY1OBB8fyPvljjVOC5BMGfObKgTzl4QPzoHfnukCK
zZSQa9dD+7tehRnhdH9B0/iQg8rA2MgXBMKnbB/XdTLM50zN8bMpe6Tt05jAHVlY
n1WT7nAJbHMUcx7dFACGbSL3cpHXvpZFy3uLftr27DrolFQFr9vzD9SyOY8/9NlN
5lvKS96wq7VsP0keqxWzHyDgOmkE9Sw8vd2g5VHzcWZm3uu//8gpKudy30pnxke2
yf4MhML3Ca9MwHeLYb9+mPv3yh5PYLFVVvyUjHKKW8C7xq9PuKQb8DqScOE/NnyJ
4EeXxxPFR/7K9wSI0X28s3wUjIKhiA36exWtgWcaDX99CRBF2RfM+w+yd2KkrMd9
TLqzVms0NSIEPtJL/NHH/UtgZicIjjorFYS+jrzNuupTpkWS+rm7fvx/DeBnRuUc
+1vY1eLBFrFieHeZvFX9L5u23KlNnQ0XfSHsqNVEWLGliOzbDLK5zy35AstM+qea
y/Hjehma8+Y6+3axw4EcDNAVixBg4Dn88FZ7IDVt1luy/gsIKEMqrhfWYv34HXo9
EbKk7P4rw15qEJ285GXWdExB4bTTO9AtutRSFIDGK6uXCIPp4bMffM2D6KpYJzgf
+8rEsZPCZh3xERkXQDOi6JXRnREoO5wYTpIHtfwO8W7iC0b223obAuD3wqoqVq6A
XE5W2dqDeoBB273bLK45FPGjBMgOv6EbS214bKR3YDGe2bRpwI3TSp3I9V7lJ0jx
jV8cexeV1v5HH6Z7tyg+BY8a9Wi09Fkv1qJ2aTWoLfgD1UdLRbvhA8Md+QmkH3r2
Um8xNu/deWxq3FDeONtgNGC8NfksSWza0pve0BhyLeuBQSJ8X750XFeolhoH0vQ/
nV8wNycoaZETegJ4ANbMieZJmBOvYLsSJn4yC11/6MJzv+EEFc+fYziCP9Z98PLw
DmWhbMVgAgkU8S6ObnHHB79+HTxphEY+UHeTmgdZ4RC9PVh2sc9SqOkilyXvdRwN
MvVAf4uUErI9SUSowuKKGlqMLJ3F3LiRc6ttpaGBUODKJV8GIw5iJrHj4qo2laWR
9E+hk7PR4hPWSXIMOR5FaKmXzHRoEZWXpJp3uLT4QBakBy8IC+hbK8KrLaE/xL3n
RM9EmPodJsHsEExtTeNAFyTCFlUWLaOEuIj16fawp/NSzHfrf8lCL9SMKTOpZdE9
z6FDCyhZ6iSKG33u4qsRTrH7SnqSpobnTiTJ8GaVwxRaK8dUlyvmGoO5w30Z2T6w
lNtLALxk8vKgYeQup372EipcMmSGTOCnFUjukZ+3Aq0SHNfFTkvyHD7bVleDk33i
EdSOkdRvAj2AjnIMmowYf69i0SRZpORj7czlFcve0FTo5KxIqTGMvh4DfGlYqKMa
9Q92zQJ4IWYupCV5DTXHX6+8LT+/qVIx2Ed0lNTJKgTwI+4yogwwZPVwoV6vIOpe
a0llq+D13KpUM4BaJvH4FvgItibUe+s55z6eabKBhKBcsuqklUch6B7TRyPOB7bY
mzQoGKMxJ7WeHs6aozBwFrzflcNhRY3tOsZMF+VrnwoR8FMnL8E3cfMij1xVQVh3
cAVZ0fKKBhVPHocgi639/pZbhhpcytym9SiKaboYJDxfLCPq/LB49e1tcmYm2XOL
9l27BecB2gc4VcaPOdzMDRZUmRUYFSM+lbEqznRmIBFqF8i+pbGOazvdeAy3/Nb0
Vn8hITLBqQO5IUKoma9TTZW9kTAEJjFPbDcaDGW/55q5M9aKzN242D9B2Z97aSwB
LrcSokL+0vXK3EKMBT5AcQ3sUhihbyfn/5ZM7qG1aDF35DWY5t4rFQ6lluALTADH
ZdlYmfvAtKvvyFLdvUlghs08UBjfAi0qBAZpo25/lg8XrzECuExC6ME3YrxBrBLy
GFOPhvNZkBsMN1Rh98ewe+ho7t3zwl+47IqFKsEDxc/fQJoFb6y7ZI+zMmOE7j1W
DXSWwSnqjwhbh8KVh62G0dwktVkufkpJHSo3Af1/eol6IEkBnZv/CQ3uyib1UvL+
iHrJBEzUxSM9XvhirUnvePLSTz8kBsZXok0GYmzIzTBDI0Ul2HLxv9j01xViNqFp
WCiTdXQF8poQ5WRjAt0z0pH1Efc6S/De8cnqwMFlzh/y2WyKR3kmldW/ObwXPJeg
Iv28iphnCb8GSVS4TVH6h9Xl+8ktfdF2jYun9Yj5J9M3HTggxR0CqKiphjJWjCa7
l0pgXqKqHzLDRDR0XgNKcu8/YFXtmDMmBJxD9g9lTxHBTU5Pbaadzkrh4nX7KUmi
IWj60APfvo/y/OHldMcILt1ovG2YF/MRAINhVBSpEZdTDI65Ef++kUMHjeozfJnb
aCAwZhH7ikSaqDZwy2/JU7VD+C+34qY6hBTmppiC0pnbwDCpTpSDCLEceJZil54j
8sL31cak4DC/DLPEjI5h7xHEOudOlznavYH86t86PCsVWVTcLRxd8RzWVQDy2QYP
IiRS6VlpWQjeNxzwwR8kZF+pBCeKolF6I4ket6U6VnONp0vMSWhodNfPRjQl2oBT
AyAWD0wD19lf/h3tYbPp6SAbt2Dr3BdMtctAqDowJfOU5eYgb4GgBr2/rccZnKwh
Kh87KpUS58ZMjmO0dQsEMhA0XCXLOkvB4N/uszE1pNnaZdVcdmedLQvNV81I6jNr
ykW1c7ibq1FvKAGqM9zzZQL3MC8I+cELLRtaU7pF+LQ32+LTYP5K+uoNBnM2uGnu
VQb3fXqE9fR8HjaUpZgXoKRL0oku6FoMzy+FcpNJbj+itT2y9ljjSPe1fpOxi4mi
Y4KdtsxMLpAzcieUOSwHwVsH6JZbmE7smHl43qD693uP612AJrLFgj8uzo2nS/j3
2gouCcfqW1OSM31yc1MJYJ6mw1VkzN0nbLDyrmlkTF1oVgpu1CAeqW7X39LLtOzy
xjQdYyHRZnHzmB+W+HfDSilmPoPygcWJNxuZzUYISz8d9yoIwoCREnQ66csAsuMr
FaZd/HrbQ86szNxftqMG2RDzdXrZqSVSv7+ItFEB6R6KxdmfEOLJ6yqOcul/uBfJ
Ex9h2uLYnHILUZjzJtKl93dBiAJC/W1wd1IadrfCyyZ5ZkYESyXE3ZDUVFxowj/4
9xNpPL+Px+bxf8aHqYMXYoG48w4t1Gn51V5bHVkrkWoO+8aRFoDYa6qqW4zK6s2J
2csJGhdw4M8CHFROTeZvHpKBQT93bXRS6nYQ/YgRElaFUuL9PiFZ/Qlkuj5Qx7F/
60QcJjzOz0GFigcDsuoZCLAul/Z2mZRjxAz3tUeHV4xJqAqWYsN5hHJeBXFyEO5c
QjqZjmgaCiPwTy9vE9xJ6CxMUy9mmBHmNwJ9y3HDFoILM0zgyfgvZm479Fq2CH1O
orsRJREI+fOTIBqJj/7G2S9AEx1griVy9HKKGqyRIacaxfIzIKxY0Uk9OUVbVqUS
HN5mY6jHSSEGDC8zYSBzp8s2/9pIvH8xDGNqwXRggOZ+MFL6Sym4sVe61ERe2fLC
1czE6pMZT/jL+3NbhIHo/q+yakR+IQDik93fguSUTuuhd/04AYVcngciDTofGOcs
IZ6QvQ9jo91AM+Q5vN1JdRXp9PdKp18jVzSCCrdPbS0cQesDUBD7z6iFPMFFaEd7
AQTr5e1eDBRvtU2N9HqxOIMvcrVTibvwFkohmO3rssst1q/UkqB85KAdG65XNDLt
Ez0yPciD/YoGMmjrKhmSXayMlHqTslLULAyWhPeue1fCWH46gfR4Hv3n+LVAcXe1
5jQWe6V6z8wP2f3QNcrbh7R3NadrCQIFgm1PGflLONQeZIWPXt3xmtciYA1A1pK+
Yq97c7HExksliCCWeQglDUSv2YKVAdti7feArRfZZrRh0NZZwXBQlZ413/tbVXcO
ofOVZQe/eND4wflgwMf0zzjRm/sbOkUMVf94d3kY39HAuc0cCexkKRO6lFozuUnY
Nw7bXgloLZlC4liHFEIwY2pi+8EJYvtAoFFTJoXXfmTUNbx7TuVVZt1K+dBbD3Yy
Q6cGH3GDmzqjTf9kCEp3BJ3zvNug7UDt+F5nWlREM9FAza4mOiZPTB5j1HHnyzwu
k8PDGuEeaPh39jKqDcrBadgy5CTGjx7Z0abjaLEQT9XL5ylxCnPOoctFHCHD+Qrw
jlGlASJSrFqYpFcS9xemW+zHETShwXfnDfcXe+0v8jk0cYS5PQqT06lYxP5K9mLq
0c4Crk6+eOUEij+GtcFOrxe8FGd/CcwOrnY4KEVpyUWncmWg2aP5aIpOXOdWl2bt
1ZTmU9zXDA4GMU2p6jvLfV08atg7yWlcG2cLd/P6JoRKa4HiLWk8Qoq37FVbeJK4
N8zij/nh/aS5/orOBNCHlOb9qOam0V+nHa/48oVXbXfL7TdHFXoTEfA7/hKZsO2B
aXNUxG0mAxbFudqnR37DY/kQRAXgUgtW8EI3nyZW41c7I3CakXCtRG1RL4ep4V36
+PWq9nCWtENiK4vS5Bq6LkSw4wDmscfCXCkQ5BZfKV5eu3UOF4bBfc+a45Fyr1et
H6crmAn4wUTwHCKlplpnCmlN0yoJHgFUzPGZZX1kHwkzrSFo7nbTfVBY/jQjO9L7
9/dhoxBeVPXcxjHEkhBbyw+EOU07ZOH4d7W00huHVSxchUOyCgAF9KMy3j724CkF
MtUOGosRUWWeyPX21trniMLBgaHI42ym+EHjVSKJTq+uXCt/KyI4+1u8jgPv5Jjj
6uF+t6PXXqngoUDHHTDuec3DLNSS9zXVNhGAIE+H4ZEnv21VlMubc8UluvSDGcKH
l0SQ8EaXTGEIsNPqq7Zrc9fVqVPpsMmBpWQgFZOijbUTii1WxR6Z12bfKf2OF75t
LAq5oMgVZSByuzdlPRUnIta3weHjYbPF7d/5MKtj8n3YooqShEOiUDhpc3Aln+le
VtRvCjCb87M6AdDlYdQ7LLz617ygEOdUzCCydDybqheJaWq1NQg058ACMIak1hBJ
oBr4xSrzOrU98g+3B8neEsrvuRxjWhrbJrNMuryCjzu6Tlk4lX5qHEA6ET4jV+u1
gRq7eK+ySISbu0+DTttH5V/UNzn5ArRCfUw7kUn9KQnyWCrdpfJtS2VJk7tynVo3
+/C7V069mjF81lRB1zAP1euRdf1lG2sZSBkWNLlCXPHifRVVeZYkbFqGrNBOlNaj
kgzzTI6CDEmDbVAFwFS79QqZSwbtiudS5EBLJ+PLILu1m/7XpbTX6pzXGIGkDEbA
XpZAOiyG+Xe0TCvwYjC9nVgIiDPC/jKHUDoOrqH7noZVXhq9QAXx4gZSkC5ScmyK
NhWr21S6w37cL7ldM++M0nJnEGS9/GSoTuMvHplObhGdP8C7XY0puwiNua5LNq6e
mTNXRUCqMgqoE1oApoDRrPgHQnmwskSaR06uydUb6m96k5VYcEd+Ws0Ury7UcGvh
KXtSfWjpmXkKGmPp2hKBkf7sLjxx7/jsUXUteGtTT3QtB5FE+TI0GAD6+2bmHB36
20gtunJ8KH06tocb2qHtqZyU40rHZLJLuWng3ktxlaZ0VlsYuBmR9ijefmKcF+A+
tp15BSWWK7OVzfX1bdIZvqiBEA9PHl7zBAslxgKA9+7JJdcKVeJbJQOQUQDEh3yl
4fQDYMnVBtZihUaTPLAega8NvAO5posKKCNbgmLQQojz9i3OrMYRKJFntoNcWoP0
42JfYJuBD9PPwyAqPqPevz09JmrhUOUuZhrpalo2+2vTccogalk67h6RSO7H/6UR
D/aKA+8xSiDFS+KnEfY8YQVoLSohYqjBFvEcze/Y15Gsv5b5xMswEzLycObEo6SJ
x7w22Cu84KbeoJiqueUZHh9ZwnwyfbOp/Iu8HsGgkvuwBPIFG4lh4HHqbowz+/rs
5FBFWINbbW/NIc3zpmtRokylNXAs2j4wyVzl5uf0LHEfa0+LsyUlGWeSMP9X1HZ9
WQqpCABR4YscwSZRh2Jx7Tu04cy0SyPMoiuA75HNHY3qkE3KH1Eqf8LpjgCO19rW
WZaPssXZI+5VI7UJJDP+bWxlZ0RCS2Xiv94NIXgJNvo7uektlXjWOtMliQKo9uo5
hpDA8TyLwUJ+6SOujYDAyjZoAigwev1Tl2uvmywqBACxjO8PKOJZwjVnCZWCCLmR
CQi5J+aK+zE0reZAIiGrK4L+JvP/zLFujySPcqCQ45YUX9OMT1vnjoE/eGcCXaKT
X7QAtr8sH4VXXEX8x3/sv67A79bSpDQnXqq8dkHGBins0+zG5pBIX4GPiAPAXoQ0
UiOnrvBJIqdWzV4uiAI4yC+WH31J2Or0q/BmFQkRmTgxEkjCRfEWDhZq0Qv/ZxPL
ggNLxZIajkTsihg04untjiM7uX+uqReCv4mo2dTOPHas15jmBX2y5cqqQQqBWlWM
P+XUbgavsUdClO5FL+Ez7ozVp6RK4WzN8xRrJBZxZ2pV/Iqj2IISqP9p2vb9c+ef
0YpyckubHKlYOOCNADFom7plh0mFBaTAU2pAany5wEykY51qbx/5FnPVj2b2+6T2
Ui0FNqZ8eElZQPuq8kEdp8TCvpXDf8+lE0jdrYLG7AD9I4rZKDpAd2IIfFbKg5wh
QgAvs0dA8psP5GRKSlspzKRMJOYXFuMfNwx7xz4fXKS8VdmWz+W/uwqALZjNlXPF
aKsVv7GpMaaxepxBwqE3JX+7zFm4afrsp5ptA+iyOxarlTY6YFnPgyGH7LP7QM67
yNPxtEmUbZ8l1qSDYge5H8DW0xTQInZZOGIOQNQl3R5u6ENskk2D0NPe+wZyHmd3
sXsouz4w7AZfx67Obicbn6Bk8TCV5WYRYkSPQBhPPPvNMOM5J/1WZIvpsIpr6FzD
c553WffxjzIukieTAHb3jHa7hMSQFbqar8mjCVney7qYD4J0w0tYQ/rEmsV6Vt2b
hVPrJTNpWyi1Gaq7mmcXHLbu9voUzd3SX02MyZbyNNCrouacDsGxqFw1GhjWxQwj
VI7SUWTNYuBm8FcAZGA5F4dgtwvx2xtyxnDWxS5tjFNoxoGS5XFVgdWzUNqvUD5E
feFmIi0NUHGsgn+mQjIDKZk1WBmpItyxOD69FBFInSeDZExDwdJoIpytTYRl7Tfd
3vKQ1vkgeZiPe5PMWJd8TywBEtuWzkjTemvRXc9MlxBt54CF3Hjz8IADiFD/sHPX
dSOmWNRN6l50VsM0PGYdN6H4ZEwLtK1BjWHKs6I9FHTzmLn0EaPVUTBxaQozW76Q
iDQM1nnwueQubB8FG5UKNv68os3X1jHn+nbH84+SixsAjtkPy/TWNM5q6pAdFcs+
fV4QtOY83Kn0v+23b/hZLNAaBReZyy68xXGyK4NmZxNC68oHwhnMYemNoU+j6y4V
rm+F1ZsWlBX2+fplg7vigiwuLuVJFWoQzVMGNbin5H9iqHgwXjEP5NbSNpnx/ujo
Tx+wDCkY3fiBtH7QwlNEu6RiYCKnLQYBILRUpdL/fc98s2HR/kEstIA6Kq0KwD8J
Ap2U3rjvXitbcg6nHQ3Kmk/jVwSCj3GHF+KJKfeotg3Po2Bf2auMtsWIIjOMY2Iz
s8nlcIrlqFu29g7Fqf5MapALtL9luIssuVdgFE6vayUZTYVSTmhTatH/cxlN5WZr
gsyDZEWnlHWJUZdL3hJj9jEiwspoQt9sNEqU8JdYcPJHcMgKbMj1BfwFUxt/sRYO
XAdRZjjcJzyE7T3SLGxrEHzpzSI0tZfAciGSEmAQqeGq6D+dH0F3Wxzz5nZYSjuw
y2gViHBr3KVtNaOa5OkC5MM3YwC4GRHCo58/NudQ+D3jwuQemftvmj2RK/sUDsvN
KJgpSiDy2q87q7GHWIQyohTxY57e4D2S0tV0Wtt8Ivf5ywXGQcx0Z/3fFdGUwyJ9
NxdLB0okx2mISqXy40y7gSicHE+Nhce/zqe0Iz7VXwjRUSI5SWtysXvmNdOAemWh
prXqIxD04h9BXsvWPodRvGJc1t/vTWm/a6xkRzbxrZH0bQAElrOf425CcQJu6aDx
MsX2A65OHvTErylIpDznrWdkmu0V5acNsFF113MGYox72M5w0DgmTJ+WYxKGp94V
qmPIsxH0uQpjy637ph86e6ikTambnbYIKlMRkRihfuWzDFh3FzAFpE1bQm4YGT7c
x4lj56uGnffWEGdyxLQRb9aj4WhER9Uvil3xAZsXJB5owyaPgjOiKQsP5W/kAf/V
lU00sfxK4hUBcX8y5ccKv/71ma6UZYLHcxHNN0XDtWskxOXZbfbC1SXL6uXS7amz
ItOFk8kU7kPrA/OoKvy3UtKwIDXxl0WLX7BcDSV0pyI1DDa8UDFOJ51GKiE0xJj+
68n2s5PNWmsqpou8xP7gNH98xxa5rlmNBMKXP8BwMHh0D0ziDfnDCt5MNZF3CK1S
MTrIRzFUUoAKBNG/PzwD0W1xxXXaXoKRHgyZYYIn6RJJfSMEKm5it0W/BcuhqDOL
JiuSOwEAovTrxy5ry/2Ut3xC/Jx70mj0kPrW3cvjS+0k15Tizx7SnilZsx3iWQsT
QPKHI8byJbd+WNJ+VEo9xrY+Rzmey7OQD9bPWVNmle9hBshutUiIp0Ry69H831ry
lNdPTp1uxWTEsNiI+LNSABsvYrLo/TGzyMDd9jo1E1AvE89Xhj4gW/alS7Y1ME2z
s6Fad4pGzt21AlxatN+m+9qCUffoYxoQ3nAMdjezk8bWWraIWPzQnQ0+yRzW0QfE
UJXIMrW0Lo1fbvz9Z5xOPDlQF8WghwXtUZSniWwf8gT2fbA4ot5gstLTGet8dItA
7ytwijse9dFdITTcGUPH0VP8WFRNSXlxYPdaPNV/0FicuExsyshClr/BktFrwSWQ
7sjPM2x01Spw8oWZfyWUP/5FxUvXUlROe0asR455LS0dbQzux11FFhXCySZ0jYUp
LBAY7D6YZ4j/ti+rUlPc5kuQX+mZSQfTONaS4y6uo2B8VMAq7mkoCyMwUbEO6InT
h/MQOkZ8/Oz3cfGVU9KnmveQZ4mbuvY4/NV1uRyydpOT9EmbT8e18bzYdqhgVVw2
5Y9wetV/+8NJuo38FQOQ/yH1PfS6PT4AyOhNSasH9WfXDpJ7rO+HGPZNtv7ZMPik
gCbZbhnq1wK/1uAyeM4XacMXuisAeRSmUqsXWWZAnRJJVo48x2OtfqmjqHNGyPc3
faEfpeuM3dmevdRmspmbdFbeWOE09rG0FnFITboeSlx4KLp4ccbZipOmboixqswF
jMt3kLeFs7bHjUKBmBlhfa3sV9DRoU0+tVQm9WjJMmWAawbiNXAwFc9THiLFQVhK
h78G3lkF2a1fnT3yQ2TSvQTaBppPnb9YzWFIpOZXCNO02CrBGzJwGPtmZRg37IHd
dC/CDQLhADE3iN1LFoDIOeSK+osmLx7NLb8QSDTVZn1OvwdnShuqqyj7pma3/rHl
k+UAfO4F/o2U9Ba6kfN9BtVQwNkRpIhddtwG8xx+SEfW+VDB0yxxEuwV6eEZ32vN
YnWpDa7QjaiZTeJY5q4KHZzwlVx2ylL7jd0kxkK5gmxTMypXwf6BgKpiuHCCi7Eg
yBbrbmzPk2+/FaJDgdY2Ch7Mj02AGzyKDOYLzIFJusNk9JNPKn2vam3Oae97Sfzp
igD33XtQDRr79nYkrATx8R8KcUIU8okvNN2cgIYjW//YfZnVCGgPNLy5fGnzWFu7
GWR8GZ0jokmyZ0ei4vgTdAKCfAanZaZYcGbDAent07B8ufVChSEXQUZ2wypYKeiw
lOusBSBgZhkvc4c3dY9AHYcOxB1pWUD3YVUctGE89gGX71zlLqwTe4BOFA6RaKq8
Mhw8Vnv+tT7/J1BEWM+zS1vcQaN9TcjMFj35ce2DdDrf8mvYo2vUjkairRRrgTGx
zWHIJiOivX5VrRdQcyacUjwlPPpwMkDkwAoXe0IzPWywa7ITLxWD0Dhut9DEzXgj
QHu/CqHhpdAIQWjyq/mt7OiR8oBi1mV5ORkbEOIWGWzoOvbZ5hEF7XN7we3l7KKw
ayNZGZjsC5/EL4XNXsZgVbneQVngHnGTqGl+Le5U385xa4Yhox0B3yXaG0kBMBGY
eC87mA8MArTvu4HQLajQeoS2aSfnnNZnsxTc08MWsn6S//ER1j4BRjW/eQL4xoNO
VC80ZeWSK1kaudYH+w+g5G7Ay7BfP/eAuHRNBSNSw6lp6xWdMDOF1EHUlVWeidk5
cBs71Rq3edQUaY4yiNcOws5v6mU/WkyZItviPod07uwVz4S9Gw2RIcDQ5gqqxj8N
FByxq5+lM+5gWam9ZLCz1+1/bSGd9RdLSTitLKlFnWJB8W2vGzC1XOwq5FT/Mc65
f8PhgsQEBOPCXQxoznqSnBgw06W0mGf0GZbWP7mmrQu6k5XNHw2tRwKjExYfhAza
KwFKdxfxWEQD7oIXorEjKaxCc6+4mkk6DANmIEkRl/Jb2rCLsLZ1B4TG12Pscg14
szrKpf66JZerjU4yWcHbUUI8B9WqSD+xF1ryugE3mwrZ1xIUyfqbLXScK+mAb2X4
C+ocqFqydw4kFbs+N5p7BIpFRDokqDGLtKRm3dPya2vTsOBQq5xWOyy8/vR0hY5d
vpdxOPfxa/SMcobUq0BKk8WULm+qfPHbvvbnsNUVlh8MycRHkVxZphM3jve6/+iN
bBgcdlVZY61h27JbMVQl4F5vukSSXcJ4on66/Pi55hvNNjWnZpK4xIS6gggz7I0A
6a0jgR3bqyfgIxDVqdxdlJOA7PYssHSkqRnKMjpzI5YZeBBZI8LxwmRD8gl6kjBX
/uoEVPysQ95bf8ZYXajDIOfue+r8ssyeAY9Yx9VOA37pJ4Uuq0T0jtjF6rza4laO
0ks4AZ5RO0bjeu9BMFtKl/8mRkIMIlWyWPEfAM00dT4OHOyA/BoTXHPXxdKyq8JA
qAg9+EOoa2aMpsIVXmXp5bAXDXYZW1VUcCti1cDUabFJOCNWWDRo3cG/asTJRYjT
syvr0BUUCDM8xuZQDZJc32S8d/JPndvlkLJS4cMl+EN+zQWM8ICMbTJZvU0WfRqf
WeXABD8ZCQbBt42iFDLpXDPkgPC+tC6Bx4IkypGdmKlzTdtIkHxJV1hYZy1Woyg+
SRWKqUQ++BI3QWTkzvmD6Y5+Aq3WDjjmInBBNss8TldONY+macYQtz+iYZD7t8sb
H7wNxaMWnrHbINAFX7Cqvf1Uxu2pOtGFKz3MECuqrAhkn6gmVfdaW5EYpraXgJlL
4+Wo3OUgTu/rrvL6CNmSnwA2G99TPn44eGsDjSyBEUbhcmFTXsEW38hOi3AUXk1Y
JemiuC9mXYsE3qRUP65/uHdPmHOeS/OYaBvPPN0Yiuko/r56QE4ybPgQl912PhAH
EdiE0Wsf1mqzuvV1dfah14GJrROCmg4zXLwsEfF1WD8rP1GOr6SYdseDxpMtBPAl
IkqdElRA/qcO12q1I9ynhlG77BT01Yxv3WHq5+R4eQrDAYFnNA4JTec9O0kFcOZ4
L+HpGydYEPYTDh+pnjpdG0KWjCK1KFEQ+DDu86Xmk55w5QC/oCPsa8KTVLlrhIhr
M2P/CSLC3tXnu4GMf4EmpyFrrwoFAv+2SihGrlXfNeuh14V8L0BfGKmx82NOF1gA
Jm8lDOc85YRnD/QI06xKQCdhAJvTUelPcECL2ukTdt+VxJmnG0ybG6sgKGXl7+7c
PMdO+6H8xDg0a4cYUMkjKmwqJt0Vwcx1YIlfJwMdfkUYudV0IyGX+7icCegdlDHa
uU0yhnaEUvXeyop7Jznq2SGXmxQWNOM0fc56pFHDYBt9KIKmFFpGXisa6Ymqn2cw
+5BsQYL917i5yptIDQ1KYgjYWqZDL8ta78w+Vniu1FM6ZTEiTHQqKH3+ie6H5RcO
RWn8gJtxUfMAoInVWdt6F35rEz7J4KEg6uZxnikbugUejfn4DfvatXRm/ZQSKFdi
Yt8/CsXe3uosj8RHryB9oNJAGcmlBCMn18QZQgWV5GUW35W4zpp4uvIpgejKpev1
1zdcVMl9f+TAtq8LC/6xwC8m7xD0qATq6oNrhIc4rxLuUI/k4LQFHEcQpiQZbGDD
w3rNrL7d4OpWzcYDzLWWQbgJCzt2ohzUUwv4MkiPajFo0OHUOfrVhl3wPuBJsQ9O
IJ8yfxjhk8sWrD5Waw+Ua678TLAF7B+veFFt6REpFpYIhqby1zDrf2axmF4tnR7a
cd2W/bjm1hJN/+AH4Fw3PvPIUPmnpboo9LiDB5ADFlFLBVdM+mmjTSIpKksn0Bxn
6u7fqZh4XhWjjJBDECG0m5sppTrE83iphwQjTaYT8EHNXZKrKMfJvEs/gjaw0LEv
v1+zK2o0epe7/RhZkseqyGktSdQ+wJjT7OVgw+2usM0/SY1CZ4t+Evsqpy+Ki7Dm
piBLK7TrsVgU+W/+ANb5AwZ4GTeNN0rCR9kLh5nG/TKKjtJivOTJy5DMlb5UkD6l
sn6lTQwmLtGV4rt+dn6Ah+RIz9G2Pl2b7GZrPaic83cemfbNe7/eEPwtQnR4Pwbe
MABR6gUs8j57sVE0DX6s/Smc750pfFFJkXWMqnRHO62NMr6+3nql2tWiL9jHUyqc
VTeSNepDm8gFsfWkE5rDQsj+sPEly/4gUQWmIpRwJ+D+pKqQ+j/zfgf9vaVrapRY
IhKeJOcbZTaVFTVxPqtMAY5iuisGyqGVzUF9Gde3Y0MsapIEMfFj3Hf7MyfVkD7B
q2+MtaSRXTF4oC7mWK6M72W5E/Y3O0FRan9lXFYNl5Yyx/WQh+5abLQ+uBc4wIha
NSu6/UiBzrB72KtEd6Rg9xp1OMyVHbc+Fq+rvELpUSS5whydAyPARERV59ASXZ5W
/YX2/6ax6XKjUoYd6VkEi1TpcgNEzHutouZBl5DpCB7l7EMvy6/MG9vydB9NYm8B
rvaueZjaOBuZgNYyN3USERrC4cOn6gxLAhbJ53KY9kstluyt2U5eVYEsKZKDF9MF
9XsqNclO2r5h/Z2Xbhf8bWCCV1rsjaILrV+LgHbeLO18M024R+F4qbet9rBAWAL1
p/7/O1jGFJm0abMmRBWqi92XtHE2vN4S2NHe5RRoBk5Bu+I9K2jRjtlg1+olHkpN
4mXDyk1DRq+Nl5uh2rvLDyA/Y2S84ieZGj6HlbMYhKa83DrYHaemCM2edvai3mLh
X+4RHXwk2aZS24KLoplo1gQ8k8jNI4SghyEMub9I6VOK77UlExYictQTcdCAXFNx
Jhtazn5F444l9bUl5ZsqKezPNdpr2ral+01TM9Xh+oTdsH5nA/ODy/e0pvXpe8pJ
05wDhuzqkrOtLIlVEsTEYySL3vWL/lABiiejDgE++xQBUZDdkURmGb0sAyZ/taL0
7soboxVGtgG/6iGLR/heCDQYeArriOzthnRbca+UhNMBBwChyROoV6JDoAengb6Q
mmdVSS5aZ7CN0CkfblMjgJoyP8Y34etOlKntm9CgNmge63ZfE7LB+8w1sZUyCpba
ioZzsOtG2BmKM6khiqFLoiB4GJTAXMzYHI0qAewDosQiimMq9AqM9IPo0zzdPLGk
JiCNR15+b+0XQru5FnGLZDLwcZJ/N4B3sYH9W4sMi8pL+cs5SnRwEBG2HJYZ8k1m
bQGOiv4EnbgX1qElwkyfzZSjcboz4+g+LDYEoUUTqRWETtoQzMcc8R6lKdtzpfdu
O5nJLmzvK1uGpicw980fWc7G3vcVoF242pdzxkww80lqKiiOpJi1Q7Wh56npyktf
XFybbBHo639I4imGxvggUyOAeEPxVsvVBvEPZOdu/nvhnwuL7yP5gdTBONDegXJJ
sk6GuapTydpkuZD8kG01C9aLcei9/ACD3gIWXwmFiS0r7PHalZu2hTlscP51kISe
vkErvr9Tvzd6ccbv33O8+kWEwUMaBwC5RwbBOtM5roeR430ua/sDQR/nJSUPG2Qo
ukm8XeocTCzsEYZtnlDqe95HbnRWbcXjzQcf1UMH+2hlS/PbNK5uNHi6Y5ZYDuDC
5lv+NJzCZymlTXftmHkV+rTjptiMEiv07olSi5JU6ouGtmlOPzIfR5uZ+MeQKFfB
YnTf8+P2q4+85XMd+j34O/5NaYSULEwFNOJ/jyPd5kpOpot8EgcBG6L00ehSrADp
zxIJtV7uESW7lEKnNXDQiyXtCSsxACPS+eJOiTWUInwzHVpgYg7wU9W3Sq8i+Abp
wn/FwQZCK5OITjkwvMphz47n8Jnp1zcSCQTWhHT9s+FjBeIcKBAgV79BZbdJR6El
au7Phol754nspk0mF6IM6ZSQHpsROICKbiU9B70ENzG3yzEdjKfrH020INIgKVWu
fNrgy7NYROkOAHXfblDy2Dzk0Ag4hDhoscNu7ZXOSDG3T8YgRqUzon9Tieazp2AO
CpOBUmKZN6c61LVjrhyAvNjl3N28rB9it5vXKCpWbr5Bj9fL9etb0H6kAlXvFGvg
SVqEpPg8Q6d0zEHh2NHvhthQntm7DNdAi19+dwNzzx/ieLs4YtFMCD4XlQrylKhz
a4iG9rRktvISR9DZAGLjSZ9564gQ87OjY59xIzQJcJdzjXD/j6B4c8s8cy6jrUzL
QmEvff+GUz+tdJ1eE5a5wsENytI+b6Vsvd7qI+vDXNrBOLRWt1p3rr5K3ck2G7uN
hi//OnbOHE6M7rmDBNyGBzuVT1LPDLSjUckihV+JWB1fbDasf1J0W3ZZt8WB6leU
dadiP5q+Pzc4RIaMIWYrCvLNzrDTbUoUm20wHeJYMPmSmlFG6m29jugGM3fveM0r
Crh/Ky0kePGDwTfA2mc+8gIeKfI6K7yCy2W5ay3UY9Wl1xiyBz2WXTn0SbnS1hch
N6iqg34mv1GAPRjI7Y+L9OAhMDtcEeeY5zYPx5YVt5YaTa2LBtLHbZUjZ+9wJZbx
Ed2xVLb/BUoecdvKTv00aciEmOJIwG26JrZKuLlsrxJdWjI3UDvmHxrIjfHvy2Vd
PrZ5qDo5dNGnuNlwmh5QYdq7NGS2euMz1Fdkc2Fn1BTiJWQRMB6yIkcnuGAAG2VS
PrgwkLQtjHYd6AQ2bWpQxFQj2bES0L8JKjbYeOIwjbMPRiBcf/YrpR/X5MfcRrbq
FnkXNFo1tdVVsYfYP4p7McuqxZEu5i0EBejpxuLmSE5jQokdj5Xq7uD1QlwzfBGC
HFXrs0e0ybPy1q/dBTEDr6F7EcvuRqhoWVyaItzYlUI99JfGwN/etJ5YkGpor2ab
NSkMDqbNIJlXTLO5ez/4KFLzAYexvg2gehuhFeIUBhYv0sRd5Ek3Wq7GAJMnga4s
qia8PdGWH1mBJcyl/PMnUEbOQlXhe5IKzS0e6smSM3dIebXNjdQPW6AclAPCr4tc
lohBU+K7wE5CIlXBM+0M5tHSYzlHt6P3MPJ6r/JawNxoDqUBVes/rVLlvWBmpGcW
BdqL71gI++U7FBfPx9DvitDh41x6aUgQDW9OdaGXf5c0rRIZtytsnXrx+sN8AFXz
R8Q2WpIiuy3Z1ZsORoXKuVvYdXx9XSkbze1Mc3lFI5n8Qh1nrZn4iy+hqQjUOblm
pBjlQpJp8cHzgtDqN8IiBNaDxJwL9py5ZyR9wf2oGGioEUI7wFHWghGFYl3OZ9Lv
tds19CdAMKk3I5z9ynC9rGDOFL3edKQdO9OJv7mT8QQ=
`pragma protect end_protected
