// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:53 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
VdwUyvCYrumuxccwQz5bcC2qcBLVGtATnCeSg3UZk/vtZTrytp2kd6ngIhXlgk3B
pNAMmjJYm2oHRQdmCiAUZrq0TdfI+Cfqp67zg+7aQ8Ut/LGrNPci0zYDfLYOKz/7
AlhEZuCvxuKB7hQS96rBlQ7DyXHE7kohBpTQ4HQmAOU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2976)
sW49rRvP3H3MwcImd60XLBKgZNQlqHmK4x/aijaggrHMw6T2HTQrzmPk9rq9q6EO
EacOVPndkK+miKeTSVIhN+mghmV8Rj5XSoipEd8zMuhDcNoUh8OmWDAEles/JxPm
BnA0e4typjD1/oGIuEYBlpekxTbG+bdg+awNiKuoPMzH8WN9MxkvCLMq5mLE69mE
1ao7fTCWV51B1GGVIxr3QZ7NKVJaAUfd2gqpr70ZkymyKcs2kuoZlOxLGivxlHP0
V1qHnezDJIoI8dSM5O5oKI6fHfNa5SOtjJuBEGaKUKo5HoCwFq2Gm3faOzo+cjSK
P11SXrgHH3FZJZloVb2aerLnEqN9BX33KE/nd4tB2ehaNBIxgTN1fSbE053LCO6N
y8PV72Yn3kBB+hnofaASFC+tcIcA5Hw9Tcg+pLlGASvt/r/GnvZ0bzo9kpsiFPOX
4bjjxAyK2UTRcnbx0uW1aVkmvhZTIL0UiGPuObEAr5A4L5khlATMXFcFyKtUw3WF
x3uUxGf+ZxRybl9V4zBgRxHIad6aS/SWWeM+j/6h6kKF6oh+Hqg5Ym7YNsu1923s
D3znwrtNWrLJsgyaxd1wn3YGZobsdrIRWo7BKAkE5LLMk7Por6MeSUesj0q1qs0S
uEuJkKZDZZEdeRXb2Iki9tgNFHUL1xiLqMkvaeI/CSBPjHMkjwBvkdSjEF8QHd6J
vkn4N6Qw3zeC9PECPSnsikbiy+S8d6NWgFToQZdjLGCER9VUABkRx0CeaICBAq9a
kbVoZf6la3n/BZjqxog5yMGgILZJcDlC2PnBAKRXXgy1/Ukh5KZHXCSApCnaVMhk
+OZGvuS2k/YA7NB46ZMrtVcFlgtrHzWKKSRPLhhwWffg0ct5eeJIUmD+cfrSmOsC
GnJlur6Zsk4bC3l3ySXwpoOf1y5spborTW5tqKvqaISD4zLkSImYf9rlUEhYrEbq
iOTug4B+FcR7CzRaWoWXpLa3w3txP30rpNwckxoS5RndkdFTYwPWv8UAdwymy3bd
vUY8qClkMijLy4NxdvoBxMKc/Df/QS2Ylg3Npwjcz0zad6VuESHSA1LJf4zj9EO5
XJvIi3cBHJZytjJGN8SZk8fNng/o+dT60K/RLms0GUA/1yYiAtXtQpJMLKhCbI2/
xJuFSUkIxp3quZ7Z+63E6So2TsKj4DA4Ji5IwhvlwKS7GSq8G6VitehabDqPctf+
udLg7Dm8CCEJseerJKvSMTA15vNIrEp4NeZ4Df8qkkN02nAZCKL4BYX5Rkvjaa0b
Yv+f4J2Mqt5NcoTVCkEJvwUQAVXt2XewlGWT1AEZShp1z0rVswvUAg9zN6ek6Xlo
v1TK39cxbGV195s12RNAjWqpGLHiEquMJXTdCa9N5R0Ms/y11QGZQv8JdJuH6sfL
GLvunnNjd8C/QBsdjjLINRmWjDT/SE+c4O6ue6JZ8RTqLmdqlhcBsRhulxJYu+S6
0/qX/RdM0B3HbJ7TUHlcbrT7RtaSISTZxDHIEAhwWML8vu7wD/TYyS5UbIYLALGz
10zeeerB3cbcf1F57IXPBj0doKsrk+iEC4mXc7FrQeb4TAQRp6qDYWAn8I3E7ZwG
SQ1mdaepPEybpkrYZRKAaRDgk+LELFIF3F6QlCJrtDlqxVAbQ3b2Fo4lrpN29eKm
U0s5MvtKFBq9mXuiz0ZCuGmj42OhursJO6YtSSDRt1ykVZoIoB6mksWy+P6bzM8F
fvZNf1vVmhH8r3iyUIyGLb8G1ulc960A37E73MsKo4rPltUcF3TM+3uNh5o7bYck
kVXdIhWYzkVQl8eVk7ge5UWbspIhQ+UqK70o1HQqQXD87OeDp+ptKTLAiSW5nEBa
ALjz9knlBaUywyDYF8e3joTIpUFD38ebO9/WL4CPp6lNUZ/HlAqQTA76YGclhOwG
j7M9ObbRPRSyshxzrV1X/tEnHjTJOzMEyx0dizIHC+3otXypX2Ouz/y8nvgcEsjL
QN0EYeWOnf70AcTWtc7XEEKzPgT88Ulw7P1U8HZyWuwjesxydc9X7rbYDWrjVwXh
wQx9NO/rCa7qJ2rWo5VAONvBGnqvde5r37vItBe9I8dUsyLNoFKbbD1B4Xni1xOw
K81o0UUWznY9L6sPDsP3vb+VgRWph/O0atiRTAM4PgGJTMCSIFmc6CYL9eIcL1IO
sQbnavJvapS1IOpRqmOTNkI9OdhC1ikxYqgGTWDfRyDBtbT+46XRgYc20goP1awB
4Gk0tjUctlTKX82srG/ThJ46NNV3ihfaH7GMScmxyt4uOgOs5KNSSN1k+qSwXpu9
fPNTOpi3XUUgZch0rNuJUhkqs0alRivZpyJ80RJnZrGr+399neQDqp22MzNsrkJk
Fs5XazgSR/xYe2JGT0ypPZz23uVV7OdNRKicI+oU3uCnDHKIuWGZA9/RV8vJdCzu
4RNwPMkSlL+CgaCglwe77fO7FgEc3xEDc9aYm4kn2qNLUGYoeKge5ihrQJfD70oF
yqvM47II0jZ9YuKTwf4n5fbs0gnlidHcmkF8DwLSUycFhE+RqdIBE9tRzk1l5LMy
hz5KmxjZgJE571rXgQWatQcpwOMU4Rzv6RyY/xpl8ySPK5RNNzNU0hkxYa86fYFP
MFM3TnmFHnRYXBgjwGtQdYHLEKrmHuvUirVoKBiJrJPGrBGVSv6q3wk7dvS0WUSj
3FFD/GpZQmab61vPIxHVFDmbxXqnul/DlYWpfw7xGd7d2yqS/W6NbPePsN02QHZL
S07wXIy8v6zJCLic4MAuj2huK3R/QbKC5oKDlawk1dBq9WJCpL3amyA6BJz5FhRS
ai1TG4xlDpIhUFOzzm2tl/uEo7s1cb7Mp6yZ2Vj+i6liknqjyiXY8g5IaW1qZUhz
6ybezB1VHzh097YgLSGfE2fTnWs19oVowMIRQ4ZARb3L0Q5E5Vdw/kjDG7P18zGE
i2UDD+H7cGcYfYoBeVKOWFOjFy4oqp233xTPADOkhFsurukkVzC+u7qN6ECBogwL
2WI9FEao+ypjq9PPAilCDdvoGcPmedp0g+z24IL1vpMCe7hQ7zX4spA/3eYnl98Y
ym83QiejCo87cBDAQXRwd3egrgj3Cu+lt1rLb7z1EvXVzIC+altrVExI3w8QBCHT
A40M7kCOPw5RTAR9vl0fT28dAZ+qIp2HA6YsM1FnnVMk1Y8RdLPw3LeYTqjQ+6TF
ZAEcUMR5yGaB5JlXyst/uTdK7hVv/J7GAU+V1rreRj8Y7cime2hRYcoLAJAIF6vu
K6LOTxQ5vqgm4SNUNfzPu0ZUNxIFJsikfzvLW34cL6WwitF278StWHf/M7WYc5CQ
+feeFBP/Eb9uRi3kk5K22Eq6+/vQ5jATm3rTqL6+Qlkko3R8QyZ0tjk0pCCDBC/s
C9qYoP5AFsLMtSU5SC+ivp4MXICM+YZjtnQc6Zncy2PCwY21n0iYZsfxrYmF4Vhi
pjR9Wl38SQ7OOW/qzDq/TMtKLC/UCkmdIco7WgodVANQgSl2hO/FjFieQvBQlEEP
vkoXK9Yln/xAx4c5BzEEzSNxriYiJYc3UGzZi//Ei4MrGaP8AYRudi6ndXv27+ph
5o+IWjTe1lkuH5cIEHV73X2YxXyJoZpb56oIQnvkxSfQ9tr1gIN2T9QsB8m0wOtB
w9TOOYA5Asj6IuvRbyQ4lJ7oRHPfz8V9B52aknkOghUil6K31THSETxkGsx9O510
dwMOpBgj7A4InjH3Ajvtfl8T7IKrbjZh6sLrdPuPr2CXeTNK2NQJrycz7Lkvci0y
7GtK3zd0f+wewmpKk0C6XrYghb6xWFPZ2/1lKjNjpbJrjv2nmzaFj6yQ6pDn38Hr
svMPKpJrYmPWss90yN+xNBmK30iIKvAAOr8NSqIiEx1w511tYGPJGNcATEuLtlte
z8JYaaksDJgeR7TA9yHPE+8UZ22nA+Vj8+wqYZmMgt9oxH4quJ7wmgjgAZD9dEjf
`pragma protect end_protected
