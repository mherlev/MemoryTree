// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:52 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
JRRTj+SUigxYpn7m0pXMfj1j5ZSvfH7ppqUWuj+JG81RFG9awAtjxHcXDyBa3dQs
UWbOs0xfawblXnAZ2eGbOoD2tt9WS1M0JuxRhKYviuf89Ts6PJOLfZCm0Dz9MIRj
CDfgy/dHMfqBPPVWc+Uj5sVJUeuH8OxsUudnpTvvJec=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2096)
tydfbnYCkyqt1Y7IeWCNcfq8ypmnRxbvSgRFqpmuJxJPF6tcRX+wlKxc7AVyIG2C
Os+L/88IPUIhJSqCPCVhZGmuV9RpH8hmmYFtJKvqFz5DIZz+JPl98x5yBDj2OkHo
7ztQdIhz8pUCh4WFZKikvX4iA84O0olu9YjKlv3nFtKpoH1VpX4E1CSae57hiq/8
vIjXGarjozFeqBQ2EmALjfCUjjxl9X+RFaVBFvYJgQdVyVYzfIYUNVTgGpw21LKp
Wy8TQsKhO/XLMmiIFJT/i0BqxUzUIkbW2Td8hUAcmnkWm4aaAxLEnm9JCC3vHf06
RTyPDhr0DmzbDyHS/u88BQuGuPoaPdas+T5d4vG133xbo2UlzMuJHKFUHPP+m0u8
noS3+Puqp7gTO2CphMdMIieBWscpylklIE1n2tteTiqqdYZP/c1Slgre9GGBuPSR
sRfVtVNu6+TDtDcThBQ7VBHrpqV3VHU8zGQhXTwn2600f3GK5xz+t/Z7bzaelez8
54A+wqbWJjXrnQmWv8VvgDs2kPePEkPetuthYXhSNmfAzR5/bo0rzKcka5Z4JbRz
sMva4ENgnDlR84q84vT+ivL43AmQwEyLV7QG69rSkDRSTfo1ATojF8JRO/6QWuNw
S914vh7RaJixxMPymCxeYIK8RVvmOwf1sVnkRwxhFExSR+ZlJ9hD4T2IG4Rij5uU
CYcKcr0sDjCWo7FH0ztQrjkbcffNWwYV0CXxxX6tSu9yTLbDO2/OwguigwO7rhTT
NK94P03TlFR5E0fBM85wHYgnXCqcYaDZSH/7mOQEFZNfu3U539qSnFLrDFpgaqfR
4ZLfo53eBm4Ufy4TMoIdqcRzcHLB+hmQoAv/o+fGg02b+SnxRaP45mq5UF3ktDPu
YpdVcXchM2QIyuK8441OXu0SfiDVSq5bERoiVfv782o7wb+2Gz7lmL12maZO5diy
ILC8ZCoeQfv7aMM5MHZZ08aGlLctPbqm+DLni8LrOw2jqZz2//ymszRNQOepjV+D
da6hLCangM20P/pD4oi1dEsUxgk0nfj3QxuX+IXkOUXFiVarCX/a3G+xXhdAqHGQ
Ds/YZ2Cl1Ga/Dn+xcjVQxasP+UiQ2YR9xUwLVvJkJ3b52QROo1lV9qS4BmJ7QpWS
oq2FoQieJ2FH/HXQdqxxFzWKDYhR0G21gt6G/lbkgNx8ns20aG1C5frADqytiffz
8W5/WG63SXMUygLZFMy4i5YpxNQeD0AgtP2TJD4Y3M/SfJykTZCbQ7GG9FczxnV2
WFdKFIUqc40Jrhq85/LH8mjh7FMMJC/ly+b397tnBQ9CleEXo8GmmSo9yXNOFhlF
3AYOFS0GaR6cD9/FIIhZHWjSFUzvg2vFtKscStYkOltp/VtPihlBetKA0bOC/qw+
m+qQOjnQWN58KAYMul3OD/0JENkukTG719qDnkoXtKEpZZzdhUfRxNOgti/GDVbP
xuft9IjC5i0J8uLPLc8MY8i4g2mPhZGNMYgTyPSpuyYGmPFYKyl8iZTIFpuO2NmN
bwkHLvsqsvF4eA/N92DmMMnNP446cHdrDWulXKYB9sTVtbiKI5O7lDVVXbQhQ+L8
esjF64AiK5UMybLF4QCfET0AhF/tjd6huPu4k2Vw+6if1q0GlYJTPLsqcw8hbb7O
htpjJmv/e2DWlvtgwrZMK7kMtRMs8fBaBZNQwPeH3Tuncw1V+OvoKvPzd3ENUyyF
y85odsZpf/ZUr/6GMBeKMSCbRi6B+erqmfmm0Lwhr0bNsePs3Vpz3zOC0mnup8kx
Bj8S7qEpGx0h7jMr+nAiPRf1pCUdW8jBi8ZDp+szf8+z8ozXnsnBfJT+tqUiy6gs
wubqLtyo/5N6Rqb5+mKmmkA/E2u5/M/PntEw+48OK+wfKQT/3bo4rF0fhQx/VvkN
ZAc2qNeRlLT3mTcGHtPgAZfKcnrAr3l10/w/4XSXhiUwJhDWgNAFqOi9HKAbgAtb
C3lvUVijr4LOVl8ha0ydWF2TJUa+IJJVeuZTOrXQOmV5qsaL3P708m/h0rVi0Ylc
0WZLzz0f0CTjhHIXPPbLpOcZI1YtM6vqQqmLacC8G9+ZsEstpQkNb44X7emCPjV9
BhqkimTHkGRSMOZYjN0ZYYdpB9Od50VaWHLNazGyOAJiWeSEPDsw3XDJY0arV7x9
gqm56mWZm6SkD8/gUGkRtFcsef/BEKu0vg+zO25myHCYfkZJD5xiHQml5jwn8l8V
Xo/NS8FVxAGYRpNPNWhcc1TzJ0kD/bv7FtE1e68O5bxDgBbN0jTZYmVJAfINNODV
5VQS1cwRLA+byo4x9axCbyy8Rsj2H11vfvAkDdyD5ii1BYHGPIr91jW3IaGdRDHO
sTxc9EtBVHaXcPSCy6iNQlB7+S6DNBtIpOlzreBwEJCrhVS67NPfRy+99e+8cNF5
zVTFaAd6UStwe1GSHSlpfKaU+5nybRnbbMqecmQm9XDJslCStI0MeHWoi8EP5PIO
2ncxwbebnHqoBSWW9332OFRwZ0CK3XfstHCVTTGYXBv5ZRNxyx4o1vWEWjhb27Ur
ovA65W3L6W10wr1hlAalVJdeOZ8zB9okAGBWbN9hiQ10mjt2ADNqYFh4s2uFunN2
pAasZqNFz7qrjyab/WjCPRdBlfspovsitNlI09wbaEgvDGjUpbzL8WMofZEyGbPJ
MEtiB1BBRm0uTrCnboUskzdc/nlypU4u1ri9LqiA4jRoAmd+SlHJbEFa4Gapdxhn
jEPLqzpTAGv+E4hrJ/0OFHIg81Xtg/BzjIIYh7avwxI=
`pragma protect end_protected
