// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
`pragma protect begin_protected
`pragma protect author="Altera"
`pragma protect key_keyowner="VCS"
`pragma protect key_keyname="VCS001"
`pragma protect key_method="VCS003"
`pragma protect encoding=(enctype="uuencode",bytes=200         )
`pragma protect key_block
H5?&41_SXK,<B@:O]D;,H8WR"_*O.PAKR 0@5^PZ^UE43??LV2>+M8   
H.9],>>K("'DKC0LRO3IZ>(EG[+,6N9TI6.%3S?WZ?H$15&,/"5P"W0  
H'FE7.K3P%UGJ:WUJJUSO-^=)3[=G]%/>)$AO,KY&P86 $7=#?F]@Z   
H+]LZ<J@J2WG_'C6: <%G(-42;A03#OM *&AY2ME60'R*-[]#_'TWZP  
H*341Y6_EH/C8:(IQC93D#_#<2@V/I#-+5D<&,"KA>D@0=&C2(8NY>   
`pragma protect encoding=(enctype="uuencode",bytes=24832       )
`pragma protect data_method="aes128-cbc"
`pragma protect data_block
@6:>_.7OD68[.#(,]@'S08KCZ@)56?/_$Z\P?O?'UG5T 
@FHD/N/JJM)%2WGWER*>+44OA=A C>\T?&Z]L=^DA9#4 
@&1RZ)!V(RH@IIL4I^VM.#("'!!??5:4$I \4>U[4].$ 
@6F#B'8LYL58,O+(/L'?5GIM51 M5LR1K$SL)8FTS6D$ 
@/HOLXXWT9NMF=%A=TW.?'HRX>T0?9@_\&O,VA*C>O-D 
@D)MGM.!<.P%QL!WL0G/KLL(Z_W :88$B__V;^3O9LW@ 
@X41<5(&7/I14;;-3M,\%&D-RK,Q*J%YL11HL+@['[R\ 
@9)I"P=RF@PZHG'"X2W8SCLQ%6E0:M";&!T:_,O4MCW0 
@&C>/"GU([!.NOI=13Y<,LV$L=K<";K:*_:5N@@:Q$V( 
@N7T;]:OC153]T<!P^6AR+]8@Q.#D%)2@CU9>DSDNB48 
@U_+T#4IQ-27U5D[:A;3A[@\YJ618*)?DWAV*L+&[\*@ 
@5Z:S($UBZ1<9'<9ET/[_KB$WT::<GIY";:.S6(%GZWT 
@Z?B%@PWCF0H%>-G<M.&DR=@ )572D7NTS,[.)4$E?[, 
@:^*DX,2']*'&K_2V"QBH:5WV1ZE!%(1#\(#=V,A*C^, 
@N*T ,UHNX*.TM=7EI-%(73<+[;6NW-+ML=PV<Q]PU@( 
@_V:7&/U6GVLSRR KF<JIU9JVYQ&QZ^! MC6QCBXEA(, 
@,(B_(-RS */&0WIRDX>)_GK6.):O$F$?U 2]G1&7PSD 
@V<?9IW(6*.Q<)DQ@VK8DVSM?]6!#$Y?>O:V3V=R?!!( 
@M96X?3LM*AES1PC*ZQ/Q6MT5Z<S\R@LM(K /SGCZLKT 
@KG7]>;\N:B@Z.I$J,%+WR[.9N<_'DH*:BQOP8KZ%B:4 
@+,-O$?I6'G]8WCA0MY<P20WO:["JFT'%@K7]IWC=74H 
@#O(XDWF6:D,>ET*](\4+=<'2C^/!Y",!=_55X@33:MH 
@21ZUL2)0EJGVTBVOF+*DH2B"#5&$!BW!8$_]@9&"WF$ 
@#U-FWB*IG;M3!OB-0%T/80:'TLT8R!BSS)KPI$YDF+P 
@Z%'\X3;.U-/P@G?FH8Y]N*W!,ZXB:)*"-)]P+-P:&D  
@'N2T:2CZ(R=63(W7S(2^DN+NOIZ^J1K*,M2O0QFFBUD 
@(?LPJX[Q^[54DC,V6K5 V6;I4N_T_6+=0^'Q:@7MJ?P 
@^B$\A6P=?#OA0>%/,7$WV:-7%I_AGLDW#C$1URC P6L 
@O&,0_YE[2<J6:2OQ)V'SO^_J>C3(%G!295)_5]FXX*L 
@+Q*'_6/0Q"GKP%D3-H7_#!1QEJ_A*89NS5.5]"_TZ\@ 
@[$W'J=O53DP@GO*6.2LT4GB6PFAO9T-,?7$%F4\.-Y, 
@MOP/?&"SQA>GRZ9E2)/V<*C76#QSK?^[IP'@S)_O!4, 
@/R&&Q15-)W_.+9V%+DX)S,!^4QP;].Z0917PNXZQ0-4 
@0]2O2AE49>_L7(,+697I!\T6^IB:K0A26\LHUFS_7 ( 
@J/[ORZ7C4.[S_?/G0\L"H? BBDQ7PPG7';315WT-2:\ 
@AQ"ZXJ\AJK"X'?8O;8,$\*K6B28KMD0A@^MOQRA6)OD 
@@0)S,O_JS\XCPX9ROA'?'EYA R*7>\<+KS,)+&J'/P@ 
@#L)7"YR5,*E:0O22&U-@3L S U2>[$8:V(5"2_-N;IP 
@11Q]F"=LB.):4$[FB)BB/<K&5P%D@'HH87-,S0[& .( 
@Q\LY 51M_HC6V8C6B1N2#E3_.=4]U[2COV,HZBMW=T$ 
@/44J6607SZ0*M@2!5W2,4K=/M/HR&")H"**O) 10SW\ 
@(@,D[M- ZV#+#$'M0#%?,'W8/8F#"GQ'MR(>&T8K.]L 
@9 Q]L'N3<Z_S;Q-K0#JGIWL4,!=*U@TJT)/3W#^GU.$ 
@>(NT@D75QP4T+TP(+&&VE+#W'8(RP9:]*#<+:,4.#"T 
@3A H0#.3R*>1?#^J@7'/.YCQQ(.@."<V+S-@_W)!\_D 
@$*1CCLL%;4/.8)>6Z-\QT@B*8;ZQO65G^U)< XSG[>< 
@%!WTKT><[:CR.4&[[LN;A&F,!ILSO=RBZJS:_A\0G @ 
@82BDG&H0BN8<5&!PWQ_MZCPPT%C0G'-1B[#SZA2Z97@ 
@A& 6GR5UL1NDA_VS>:ERQ;LC<DB"H<?Q6"Q[IXJW[M0 
@%;13,^$ULHQ*>BZF@,\(A_X@1D<4D0M"^&.TT@1AO3L 
@D]HEN.@JQ#HQVJ:9<FR4J,AD3I2/8)HMEX95IJH6!?@ 
@$&TX>S;<6^M![8!DU Q0L@-H_;[G7PB3"1#9_TO3S.8 
@RX0ICQJO9.9<PP]7IRZ2IZ(?:[0:G[W+[NIC_-NLBI0 
@$_K"A0S<A)E0JW]4/?9Y).Z+_9"8W".I__9G"AC?WU( 
@352R-:2Q(',Q8RJR"NU+2+-Z&3WL&WL#N>SK8:"-\:0 
@EQZE_;/ G'4UWG"@/*' ;_IDIZ?J3W9[+2E+/Z 6)U@ 
@S1$X)4^>OG[GHK?G4E[<'[4YON=TUJ#M2]JM<&?IC;T 
@'W^92;C;1$V?**,K/R6M$_<8F^4(T:_ML3H.I7N(-2H 
@3,@?VT_>$TI IG6&G#08$*SK"<1^OS^0FC@Y\KN#7$L 
@DJWJSV6!0-;W?YSRBYM; VJW;V0U$.?B@02Y"Q>IU?D 
@*ZW]!%;GV$W(%EJ(^*J9&]A4YK*^L_&V1B)$M89"%64 
@^YP6Q"=J4$U2Q$]8)8K7,OPP,6?)"_*(H( JN'H=Z*  
@ZH2!"31;*HCTQW^FU\B+!)1CH,"X\\R2)FFN *UIYP, 
@+OO*7<DSUC27WR?*RU4&XY&<NH[X&.C_K.8T<01&9@4 
@JU=#"+K?: *RE*0I%&Z<6$G&(U^7J$>8K[N8R3<3+($ 
@!6WGQ_:1O,?%5!242YY#\(DR%&KV3!'?I*=)8L,O62, 
@!03Q8Q)FJQW[8FYH3;()9O54.:E^4P)/V5%4C,UB:Y< 
@GT0K1/]'A<6/(*%M33N*$7'Q"7=&VJU$1W\;Q='WI1, 
@?6*WP">1(J3 EZ6Z28,,-4Z%2CD'7+<(TM><MCBLTLH 
@/LF?,<H$\AW'LN(B'7QE&&M29F,@XF@7EMY+F^0%ZML 
@9Z!LCY'-<1RZ3\QIL_T?)W1N3]_\A'+QF-].=A^!KH( 
@.Y7TD"HX8^RO(?=:*J 94LTS-]XG$):\2\%N8),#5%4 
@\/=C;X^)<\&CD&_@)O1]"7 FDU[M[>(TGEFX<&S?G-8 
@_W@YI!,"#6+[P:,/E?,.+#6I#TG>Q-)O#P,[H*5GTH< 
@*>>YQ,>PZDE%TP&MUP8&Q2%&DG(P@3G <7+TV.*"L-D 
@AU2N?5E&1:\#6$3^$R07_''EG['H6N'\LSHRPR1[4W< 
@5V#II5  )L+5@:GKUTC=:M0#@$C>S;GPLEB1U175H2, 
@C%R6LL<)*Q^YZHKDT[-_KL"2M-F6X[_JI'-IH5E? <, 
@.EZN:3Q 5\:Y&: ).2[)ZG86>S@N'-F+1W&[&QE"2C8 
@B]D20LE;D),Y$_3;ON8*,WQ:+3E,H-"-Q?_^A7.CB8X 
@G*=PM1BL2 0VBJ$9^\XGLWXX^UQV684V8?[E48VT$7@ 
@G7L)E^9YCY914C4;*@*#M%JR*FR,1M*_IL:@D:K@>"H 
@5ZC82L[OJ>W<X.M0#G\L&[D'IKP,'_)PY;5 !2^K=)8 
@22M5/Q?:MY,0)Z*W^H;B0)N8_M[E%)%W$[-:':695ND 
@4O.PR*OS:1"+E>6*GQG.-^EGX\98I'_/9 X=:475>WL 
@MVZZH0>'=VUJ3F, +\:Q5W=8%H1IQRFCQ0KL' 8_6"< 
@QS'Y7)%QUQKZU!G:RGXENL92P6_28U=;,7YED4/.O;< 
@;F524@W1%CJ"(AVX,Q0:$LW:U5/2+&VGK/+3KCTSB\P 
@.1.':F:3A NO3.UR:!-HH(VV*M P?1AY-_,<JE&:TBX 
@0'LY>!.T3^!&O?().4EKF>^TTP^R_M,ME;^==&31<XH 
@"H*DL3@B:UR"7T 2FLU,5:&,I\;F27]BWF"9YOFS/=, 
@TGLT?N'F54)[GE6VG1$I;7 >[5\KZ[XMJR;&3G7V7T4 
@>'FE9:@*Q$A=)?5U]G-V2!1/H ;4Q48WN:QPOIP9#%$ 
@]>ACQ%9 ,RDZ-!S+'HUN<; N44;@_LRN;) 4$16RC#< 
@Q!6^"IRP@)E,C-VHB7*X"%*(6&L4JRJ*.01Z2.M1E$0 
@PSG6[V;:C![9_;#,B7X; LV(>7#]*8=[ H"*+H!U5BT 
@FK0UC.3WOOH0U3A>E6""N? X?A$[M%@^X#!TE[=?$6@ 
@O#!:-/^@VPP9/2_:9:HAN1(3@Q6N9K-"6M"F:ZK<8F, 
@HS[YG6XSI(6?[[:6ADUEC9><YG![!UB-U!?RXFZ\]70 
@7DI!9N=MH08E*3Y0D!E9B*O-N>ZR"RO:S?97F V+$Q\ 
@\K$A%^K/4);1HV>,)P.5Q=LU1YY&_*2^<--=JV 2C[8 
@#8&:?!GGR95C#-T+ 3;JL+PZ\/6/LQE_$#D*ROVC2DL 
@B6Q<&]0I?L)P;8'X+4QR7&P=M.8E]5+($8%WJ<_*^NL 
@')YO%XY"\]_B&@#57,&M>+K0S4#!1BPRN="==C:^H5H 
@L.+)!P 3J7]1:GYV7'R5L33S6STD#B309<^@74G$SA< 
@Q+P"(/B(RH>($:C\R/3'P4$C^%?KTT#K!274\.$%2A8 
@>=Y2)WU4 MG5%1'G<76+-0DH4?/!W2"AYREKA-%>!KL 
@R=@YR3$?X%JY@ -W#O#LY$4?-,]E#2@YLN;*%7HQ3UX 
@ LRN3=8YG0@]%AY)0.#8YT,JJ7RT1\G,DM!T;G6<$6T 
@V;LV?^$QNVMQ\71Q>=*R<QS.S6^:HDV]QR >>/"2G/8 
@E!_'K7W-(O^A],3(U1R@X&(DX+BK (80VI\FF[6UM3< 
@ D& 4R/]Q?:UC\XIM(,(9MMUN5P]"G0PBD=T<[-+T]H 
@/;&]/H$N$(FN[ X7BHA7A6HYC2>_K=;)5G!D$[,MD%P 
@K#5G+FK-7@<=0 )!>=\$L$BMX>^HGV= [+E% B'^:F4 
@Q:C?JD[ L%_6[PK%'#+[X#42&]D]4;7[R,>,DN1R\[, 
@F</;*R<=Q_7+00;-T/[.M: S=L$]W%"%Z_&:Y\S)L"D 
@EO2BGY>]?.$!<X53O[P5"XUXFASGE!T(+$#[)M5E)XH 
@&F)[2NTH5>!6)FG( :!6:6U\LWA? H5)_Y5H[4T0'IT 
@AG8:ZT,X6=;6<YV36_+ZS7+&_9@R=<(,DRJ:]\%D1>  
@8:%706'1V_FO&Y30\P$2S:,&6DU7O**.Q2CQJ!C]-3< 
@RIA2M0CI.&,X6F)?/[&_5J71TE_L X"Q5O/B[+=(M)T 
@F7]5A!F3^<P0A!1XX49_T'7$&KE>BMX4UD^X84O:G,, 
@'XXTCK[2W%LN,>6$K[EO,X-!XEH#U^IWUB:42$BUO9  
@%NI%TV]0T?5'-W.7^$A][?'XJ@T\;Z;5 I[]!DH#;T$ 
@C&IP0 5E4] (LL>]"9R[FEDQ#TE%%!T%[.WYW=M(P[H 
@PDM,9?U$/JX39_=6X$?X<?G8WMX2?4\)"37++;X"QW< 
@UREGXZ],=!G@( 8<D>6639LUKIL*,ITHW]:I"RB!(7X 
@'8:Q:IU1?!STE)ML(B)=%$<B!PHP)Y))-3IJW=9B!!4 
@IWQV0@#9]FX75#-PN:?$"6K>T60D>E#Z.,5&?_6P+Q( 
@2 Q8N9OO!9 HVT: W@!;"1^NBXUVQS4H+M:56^QI<8L 
@)W;!R).TC3C$4N21+-[FEP=@AW+B;1H4RPP6[<Q;83@ 
@]>+9LM%PD,W,Q5W/6>FI,8"*7YX4N!R:\-6(3MFT[]@ 
@X[;T,[;EL2):T>FQWY,7HBI(LA,ES]J#)WBH3; -62L 
@P5LXZ+H3\'K-(;-($KCQN1] (00#)WNQ3!J-I+DWN!T 
@)Y+G@3%\BD>@D;ZY\$]>2.B/$^,O&T?\G[GNKI.HOL< 
@0:8 2%VV%NZG+SEC .RQ'3'^U9+KU:7IKIQ 1,*\<+\ 
@A3RV/HD -U4VU9%LTL!<2F62N6UV/RG[4G78Y71J0!$ 
@WZDNY"]2RXD!!C"@#CLZ1@IJB*\ 8==%E4 70\G-1%H 
@^$V/,6LJ(5*1-0&-5^$DD3%N#D5PEYB][X,;C5GY$CL 
@Z7XLU!,0N5O7QFK-84F'HHK*C$--A&C0)?8^2>_L NH 
@B77(+@<(B:\YL.C:D6G&L<B ;Q5<]]B".'.K@I1PCK( 
@24S!Z-\"!3TW9 !L_$#RX4(GG.)PJ94O!<%OI8-H>60 
@$*MZ#T",9X>HL9@;9>TTC+(M("H_H& 0NON\ 9S!]=< 
@A+W 1M:^&Z/:2H$DNA2BBPTK-A/M]JL05K6%"-<W$BX 
@)XRX 0C#S9L-(C=$]N8X7LP+%"_18P=_!\0K^MG.4/@ 
@,-,MRALL+.I<=.&\2;9,2&83A#FAO5:IWME<M&+^%R0 
@E >G$1L]RL\'UD-(HFV13WL#2?A,=KOR:J2)0(Y\I/( 
@#:'X6XY[>^#YE\2!_QI*R*N0M7.Z/5^(JMGQC5P^*&, 
@&TOVL.'&L*T(VI&'EN26R(+&#-^68X1?.L&T!UJQ^JL 
@;Y2TX<HA'.%"@K]JJF'UQU$&\T@6,M^+E)/?FEC%-7P 
@$5%H)*4UWU:/J,::\]3-=_,^MDE'HFOK0;!(V $+07< 
@=^+3S)HQ31ACAXO/N"0>*AP"?,.T26=M09",8S%%;N< 
@[CS%N1E,,"H1]T18I")MA!+\Q"%P01)>5"+M3ZG-1C< 
@*GYYX$7&KEZK673S+1HY#!PCS-4$-TX&TH;D;\A%B9\ 
@^ZP@V^Q)1X/J (MR@?7=^5K6P@)$_%R=>8HQLW>2PSX 
@,44SE%FQT+Q\3A,$4MP&?O9$!#@Q66_=(1_47JO&(O< 
@'[?2C)6=7#%P1')=CN]+4M?4] 9ZG3S?B/^(=F5IL'8 
@>]K[_ BT[[I(9>*;'0I,;[UAEF2W(X-Z6%G=IW1D#XT 
@31J1VO"2\ @$?5MZH<:&Q,T1GF^FI)W=?DTDZ"/11:$ 
@]UWB!7<]@!;]UCAQ.9LU4FE/QHZ(^M#$FQQ-;R&XM.P 
@I'+EXIQ8I[,B*&JYR!'J21'S2QQ5WZ8?:A<DGV6[F1, 
@R><[<^IH_2)0F2IUO*?=SHPD.(FW>@8TOH@DLL[*^J, 
@^59GC?DG8U' ?6H]\A_QOSF8W9EBKLS)JG=Z(LU2]UD 
@8=L?W.1FH[+62POT?!+A5W@-RK0^#*@MVW'X%?IO"2, 
@>@2>J2 E J6.420ZRI=@A9*HAE/I2'5.P45ZB.[2!DT 
@^^'5V"JR_\/=IFBEAC ,&([^\,5@<)ZQX=/*.47E8S@ 
@>1K.:UA9M! U&S6]\#0A*21@<"1DB![JZ,X#64^FU6\ 
@VPO1!RD5[#Y4&[P#[<(<;]50MI&#K?)N$FHK@@'Q*!@ 
@P/= \3(KQ'ORYTULGNJS9MIC.[E250FZ*N_+0U&*$$( 
@H6/AEL-U9?7?XJ>@VJ:GW]Z]@_H2U7Q-S/_][U^_#"@ 
@7#TSQ0']YE5:/Q&3' 9BVI#\Y-R4I?:'10K#+\2ME1T 
@GGM3DUT8QJ(]45>E,(O+"CR9S'0364?6X&7NQ!W(1.< 
@HC0&K/M"8E* GC+5)2%WKWO)Y'+$8I7"1SZC#HT?R1  
@[Y>?MU$<GBYA^:.2EZB$$.$PUR]K'T +!Z19S6K^I/< 
@>8<W)?[8T)*+%-JL!1/6:TNO_*1="=(U/HD UU5 3YD 
@"BUK>I(!RCN?,CJPGEM7:1GV?:+?OYC,U_0CEIBFJ/8 
@P70FJBI=_BER_92)\ST:J@$* 7.-2U2H%X6Q3: :N@0 
@'JF!5T<GN(5$RF;A=*ZR.2DA2T/-=**R1'ILB3LAG(H 
@-KY]-VN\%%;;:R5);3:7?AE3>2/W'R=D<D\@=5BEW[D 
@",.1B7)=_L^IHR,M5DPUUTX]7L:+*DHU@&@K;DH>Q3, 
@[,]?:9:MV$Z?'.YQ)++UA\[NR7KG0@*@Z4KY?-A4 .$ 
@ASBW8=6/7]S "CI5TR_+GDT<70./Y.F5<&E#BUN\16P 
@O&YF76H[Q]9KHU@TD)'S:O:?2%XD9L7^C);E#F#,?%  
@BXQ<\J96+F)Y'3L+,.'AA!8'003"<'*<^"1S<)C(H+H 
@ ?*-W3DCMD-C6GSB/,F,PIZN=Z)^?M(I!$^O=5J:KB< 
@QS\;II0D=<'W7L42%!^_KS:Y/3Y/"UC' ( [:XE;UNP 
@$^](15X:8?+P<>5B9_/'2H.>6UA8@7%2?FHPG)/]GPP 
@<1LK%X];1#=3DK\>Q&85PLFE=CBEU@,<$AWG>>(Z>OD 
@90Q2@,*IU0"C/A9;H5,P37Q5K#PM?6CAO&H\!_2LX/  
@F&U\,C4ZL"7'A&9*H.54X-#-_J>7<T"$W8\<G4HG4?8 
@.V@TR<LK+KDI(M3M8NAT_("0^D!O?C=R#T5[=R!0).X 
@PE!]KP9V$KKOGO1VE0?'1[H9PN67*[<JRLFFN\&=2,H 
@FS.H?8++' N0Y#]K)/ND,,VJ;L1*B \IS$-7V LPU=, 
@K!4J9%AY1>ADWM0K%""\H*SL K=1#Y<SR++M^8(UCL< 
@EXRL2 &.)9-4Y#$S+M-^>U V<69D"<M\ZNCD)77]V^$ 
@GO;7@_(2W:VBIZ3MB2QBJH3/4E$6DE>VRV9B;I@.S:H 
@7-XBQ?+ZD!_-)ES?<#Y9#4:(#3^CR*!?84X%S_'\0BH 
@^N;E!Y*+F^LV]*X:8I#231<Z8-M*C*B=T_\$6-X74QL 
@E=_?T,<3X>B)/B,FZWA%0[W.[;8S'^ (D=-AJ.R_>50 
@1Q#4R"QQ0-1Y=_Q#4W +$]FFW%77G-%I;L@74-I(!68 
@.G_TF$A*6/*"*DS0/Q]5.( I<J>"9E@."CWQ2G9L=9P 
@2_STCN^Q[\JR6R1E0TK'IT:]KE?4B.H!&CI_8%R[[P< 
@VSW8]%4TRV7R6JF7=(+#^;6UYK%'S36A%J[X4+6/PE4 
@_<9[WNLU@)ZT^NSP^Y'."]F#G[$D#<>6&7,JY!#%0]0 
@2J[MJ60)+ZYYX[/EO++V *C])>@KXF25=@1*UJ%@%P, 
@^O+A@&]^U0#]7NY;P^-E_F%<[?CG'M_[""TX:EIG2M0 
@K/A9FS>6DY<D5?A8W(PM:4^6.=&;I&-29N9XYU0<]Y( 
@I0$R_5?X54O+.7&#/F];694%:?5?"8XCQ^"KER7$M&\ 
@S.:QA<RWZ@>#R@2[: -;5 #[]#_5Y15]%*H-*B??PI4 
@X@?4P:PTMC&R8VBIW93T;I$O?A_47<J7S,<'M_4O"N( 
@E ZA*@IBUFZOP<*]G^<[9 ZSFR9O!_N7H<U&TN1F(;4 
@1&;'*D]$"+DE URHX1QHDQ7YQ W1AU8G>]UB27JBA6\ 
@)M$UP&F\C%*#SCV_CXW"0H0@)]LH@O!H]R&T@U1P[1@ 
@B6GR>2LT/=%$DP@3DA2UG!<^OQ%K#TUG@2=<1H9,2 X 
@?<M@R24/%+\T+'*.,<]UR:^S%A,Y$DK.J'*&^A%4[T@ 
@&11A*:#XAYNZ>G>@/$J;2.82F#GO@ SVFUB1# Q]63H 
@E0'.\ML#_2:VEA_GZP_R&+EA'K?A*3Y]Z9*?P?L6\Z( 
@GGFCT2M**S:\DOR!FIK#OZQ6_2-T/)N+.OU".*[Y"50 
@C>NT??4P0+$*E#2#&D \=]M4JOE9 BO]LLG=/NK=D#  
@I$G:9J"B\HA_,$^;7$Z\A8%KF*?*VFBD(\9\O='H/H( 
@@U4F!6T,C5[B&/U82*-#&R-)>R=W0.:IJ>XI8AX55&@ 
@_!@>\[%V43]KSB,IVXLEXGM^2<D'K^<ER/%,H HG-,P 
@=][XI'DX5-2-?(0++B,/W)M(+N1CRYAO/*Q?]CA+-9P 
@^]614)$L%3?WN?20J^Z/5TLP41 $[OUZM'6YT>O59:< 
@KFE1;P?R+1RRU<H%/OJ+I5&= F(\E:['7(JAPH79F@T 
@1C5-W@T?#^(=*7K7&'8:PX:VUZ-.O7?]]*S4?)XGA\H 
@6=@'S?-"-_*8XF9\9SEDDWQJ5<AI//"$J<.:72L?Q=, 
@AR?T[5Z<S51G,(*KVW T.Z\(P:PMX/9\?7@,:4D.0U4 
@>0-6]0"QZ^-UAK1<,#C"=>G=G431/?-:N3J$_&>LC&\ 
@FZ!"@IAHEE&NMY)))K@!D[6X#B#[1",4L!_5GC+@9PD 
@5.%G (;QW'C![R5+Y!ZC2O=.0!TR$^+$[D:%G4 D074 
@LJ.8!+L8<[]\"I496?T&7-BBKK4Q7^?F!IU7/TO%+C, 
@V\Y/RO?4S_L9OS39(1:4$ !X=-S8O4K_SV,&F56TGD8 
@+F]@JZ)'-UZAJ,OWYJ;^^03W%2LB$$*(,E<X?C/;Z>0 
@S&6NX5TZ;=!4%;9?+NP):,&(^C P%_[A8@J:&XPPY:  
@?!U+>8PE_-&P%@XCILX_F*%=YWW#A:&ACGKZ=%1.4XX 
@O@^OIO:,4E00\S1..]XY10BRS=Y4S(Q;I?C>=+ 0:7$ 
@3L"'1U:USBPB7<$-$L3%)_:B_S4ON5];C.ENLY%^+A8 
@J#SQ4#8X?<SL>F=N\ULQUE?/QI;<G(4#(^FP,EF%U@( 
@VAI'7(I#E8G9)$![W;)%<A]*C$'!,^_65;@I!GASL\( 
@I#FQAV^+O*&4U5KY"P6M(LLR.0?L1)ZG$F+DQC["BA, 
@,:5IVB%9K'#SJ$=+,+03Z+3+5 9M!"=)#KM,9K3ETX$ 
@-(<ULPM/G\/%UB*O>R*[S":C .C/8"V'"BAMT ,EY20 
@+6;"^K6O+%)R6;46NF]"S3P4'G]A_N, %=2B$0?-(T0 
@'M^T.8-$\);Z#'I/?.5XB*-QY">'*6 .WY.2\P('OF, 
@5EF@Z746W1C&^[ 4@#8QA%+&C(Q8[PXC1GX,T[C-BQ< 
@CJ/H'!TF",MQF3DXL;'\=M*A(Q8)V3,&W;O>0I:UHR, 
@\6SW!(!T?_K\:/%4H7':X)\/2H;0>C("%CF1N+T6%;X 
@IQ(! +-1#\F$&#(2WOP $]>&<#^5#CZW4@8>PDQ?<J8 
@5P^#V ";.SQ.[&YC[\51/<[3RF--KF+YI_)6^L'K4PX 
@GY[Y$76EUHCT@DFA;>G4M_\):D:4YW&,!*1EIXB?]A$ 
@AJ_.%2F5XP+MY@O5<SI'PMEJ,B:<NWW%H>Z+JBI31+H 
@*WW)9"D \IB;T?3_U@'4"O4*QQ4?L304QZ1:,[$ 9K8 
@]&<V CKM/"=^ B9]S^:64M0B4OM $H(W"UY":';2\KX 
@>1K2]ZKN$/S%\063.&L2<?"6;Q"$E=E 8Z_2V67+"F4 
@D=6@5\U!/3*78& <&V$D&LWZ^;/NA?HPN&V1=%_Z_5< 
@P,=T4^#;_1Q&?]^,)3PIR[BW']5%O!/9?;!PD1 EQDP 
@["I,_S(E[>F/? O/%Q<DY:NX$A-75VM-D)=5$\/!X;$ 
@@B[OX=<7YV V&*(ON5+ X-9H;_$P?O"M=(1CE%/@.TP 
@6-7F$0U9I+,;GCS9LD4W"5%NV:ED .B7-Y'*\Z<*/*X 
@"<:08.P='3%6EZU!!83P<Z#O_21<^#2N#@7%P$H)Y=4 
@3.<68[V GT9V ')7HO73W#:KVE,>7A+[)A(ZD&Z-G^8 
@,M)(U$C]LP(C7HC=Q1<4$105<^6TLT/+(Q::X_$]T^P 
@&T";\U0UD"&&;KTG&)R,+M;N3!BG@#U),QLS!=VU*C$ 
@HV957$A)DP(VZ4,UT"BI'",3N2M89\@0*+8,0S)<ZQ8 
@R1W<K53-MUAOO%IA2[E0C#N3PH2HNNDPP$,8^V%@E6$ 
@KG,ZMIYPR.F>/&1VQN%*K:2'R=L*K4'%6&*9:(]_$S8 
@-A[OH-H/^ZVMK[P7;J0WGQX([0J'VB=ZNGYX2P]O3!8 
@PXFYW".B5TWJVQ[UUR7?U2Y@S_Q/#93:2&4&JA S[K( 
@/Q@:"^_QHXYU;4O_<$-BW4@<@G^\R-G@ZR0XQ.PHE1H 
@F_QMT9-5U8DI'N#4*V9V!>MEJ'UG#XWW"@,4LU^F\_0 
@8@H=KI5 (#-572HP#.4MC1/P:@3"\&WJ<THH2-'E#]  
@8![62-!Y^S+>8"<ZP/LE[6H3KP);]XC)RIO_("+VC"4 
@C6-O&X?0W:)[F:S%*L"P <G"O22&>NVPA#1Q)*,\_'X 
@0/=9'!?7UYQ$8#B8WB/3F8O?T6-"),47I,\''"170FL 
@"RW(Z87K'%*IY_SUR2NT SLE_6KDED^'^(V;9:5!Q1\ 
@\*.O1Y\ 10,I_D+BR>.U+?Y)M:G$K0=G4J##T[R1/\( 
@54UD/*'J/E?Z#HTC89TK2H!$BQ\T37L<+*CTT'[=N@H 
@WH',NET+-P"Y_>']XS1<(SB< #^X)WIS'RRJ""V(7Q8 
@YV3.K1; 6AT?-SEQ(3O.F(T@K\VTO,_/G(TI!":\F8\ 
@,YFU'*9,;:HK#U&P/%A6DC];1>/Z0FK^KO-.E47#NU@ 
@&/5&#'F!P J\XQ> %/C%#R0>F:@97)?R@H3YIX3>^/$ 
@4#).<PIG-?@W,F7ABP2=9M*B35&EW] C4/XTUW]9IS8 
@_\..L2?XR[7EPV(M44+O7_G[TJA>QSV]B!N>6^0+<K, 
@"U9BSW Q_&PW"!WH(\\#>Y?OY?]-M\53L>55?05:!>( 
@<7[:N-X&\3YGFW '4]X>-&> O_(.O?:I*7[LH- F1Y( 
@ 65T0/P?WPXD0T6@9WP(QFH(>#TUHS0X...^M9)3C#D 
@&Q4R-ELY#@'$T//$T3=_!IO)"DTB.71!1*QOTL?]*!0 
@0?##_O@AR*H>@'XW8#J--4U?(:8[>$ 7J^:&M>?H$W, 
@9&"(0]I(A\A9B;UJ:0O:*&>#YL;M.?QP?H]EDSMS(#8 
@*V#=HV+FG]\>UC>9TH(QJJ7A.+>*N#H1B0<UM,.*G\L 
@R)B"-5IY<",HM&0,/\M\!F2-=96L1HF^=Y/BJCNL6O, 
@=(JY6->)=*;L"QCTC#P0C?5,B#:4)'5T#SJV>^NG'-< 
@ZO>.5(?5K1O<K32[SYNH<X35+!#7!=?$(=G:X2R#G-( 
@=G9:9F25URG-(\YXGF#&I3&G1JMZ7=D'8'M[1UG>_P0 
@6?,$.&"+:K?-9BJ"W4^CNR>:9AT4_:B J_=UE#'H%$H 
@?D:8H\<BD<C15'#=M*=X.V,ROB>GH.K()L)3<I2]6 , 
@H_U,'89(^;GB-%B1:0XY01RW')U=&'HOBZ2H3_-&7O8 
@*[=DJP:+F@Z8U(@UO!A_+BIT:=Q'3TDXV@VTDOW ;PP 
@_:S';@-GX8-["W/=?MCMW\AO"[D\V5NG8OVQW0>ZUJ\ 
@RW5^]%3P""*A*Y[ZW\;8PX"0T(DI#7T A2+3(8D3'W4 
@^-CN@M%NRLCV@CX92"CC3EY>Z"^KAOH<?[W'1 _K%Z4 
@*(1@"GS\-S(;(7.AR--G*/N";>/T'2TL,]T BM[P%(D 
@1RJK_1$F+Y/=8"3EV7Z30"PU)NYB.3!4Z4'@G<&8\VP 
@!1GJNDDL#]N*!TFK"'%D.V13R1GZMT9_?P# 6$6T -L 
@MRUB8#P1)EU8&"WGDDT9K[/&'@OD[WQDW)QW :;&(]T 
@. .+;5YFD9DS3^HP]<A*'/J@!O[)>%;N%3.TZI.IW;H 
@W 9^%2>%P+".+1L>'(A$IL7X/48P7F=WJUY-H5YVZ=@ 
@8&<1@)[=]"[(K=G&]GE'L(7"6*DEHP*OA">WUI:9,&0 
@>*WNG;U@23\#5\F D*UH8#&VI)[5"@3/@8MAK(1>*N8 
@!SFTFR [?2K)CS\U]1+;I+4VT.H(UC0AGI0@M9">WCX 
@0&A"]->3O359"7_R?B'+IALL<Z<#%/'[GO2=1K&9)^T 
@C9#'!&+NUK5&V<4K*??&S-@_:Z5.41F)8I&]WM$'\2\ 
@^8>1,  TAV\[N4"&QPCR59R.\JKO"'@H (LT[K2XQ;\ 
@5!'52Z2!""3SZ]G:$Z&1T_3WGF\Q6,8(O4"7W8/[DAH 
@LJBK1O]:FFX]LPGA3!V+ULL)&XVC7;E_!8,+3"8/>T8 
@3M8TV9+P/8P*MLB&*%E'>CYAWX28-FRCH'^!%I9+LY0 
@"V=S1!HMV,YZ.8;XI\7X@GB.@[NQM[]56*;-'&3M8#< 
@@$467.7=A$8.RX!7.U9?K&K=@$8PXDQ>FT#.',D.H<T 
@KI"W;!IC ?[%_#RU&V@E;+;5$:_%/ ,,*/6SN/[\=<T 
@7L*N%]T;^,YHC3-5_?5@>]^-OR:PH:5H.MSC]Q#.;_D 
@1_"6061#IO]<>/E-NVC=E,SBWKDS 2(AF@C?Y,/C+[L 
@\CR=W0T!F^0[[1IGD=(Y_(0\#H0(2%U,=8.32L_8E)\ 
@[6QK5$KQYHAVVK!25W-7]-\T![7@[JN;$2-F"#CK/Z8 
@1'R)XNZ=F,O3E%#G1G.%<B=/C-C-HI)!U4K[>U>*I9\ 
@](09U&S)[ .5IWE<?FP)%R& OT!W6[.4<+#7><+\B'T 
@(='E87W_9QJRT\D/0YR??Y!A^(@=]H95G3)KM-/A.J\ 
@2W -F\VN>D*)VI$%5E-0SZ''^/M.;_0>]W29UO87[K$ 
@4><SAB'%/#E? 4:D&$V;YL.9>N0I+*H)::T:/&#C8.0 
@H&PX*(&_XU%K<;<"&%>P62U&/,M!40$&O?2OAM\!E&\ 
@P#&PLPU&(<[UXF[;0TG\%OQ@_SK+"#D3>2-XMR9&F T 
@O< 1_PK':7BTH& XV.%"11!>.Q(*[;6&@<@E[#QT_;@ 
@(;;FO_$3A81*&#>CUXD03P#]FJTU!,41$N<IWFHC><0 
@^< HH95QR]B+DB8O'*AJWL?3@2)WOF:2W.:<>/,998@ 
@Y#=(#R$<SA$ 81<8!QZL!6$=C9!;X81W!Z,RM\RQ&@H 
@Q&7\!Y9I'.$L.IW5(18;.3!&H)NZ&'T8'GU:GU3\+@D 
@X[UME?@$A1'XPWE7!C]5O;L>.OY[RNK(6(]4"9RII2@ 
@:F,\@G&I]()=B?4$8W2![VF"B*K TC$5+5%CQ\#>NA4 
@QL;VG,Z4^,-LP19V=O3-X5O%(GJ%_6ND>&#F)J.@M?  
@AXG.L$K3?YPFIMZ5YS+PQK' ;1-UW[E]^0;6')HT%6X 
@2FYMA&"AZ-_H#Y6C+(E*A0 ]K%,"0T+ GX;AMTQW!&L 
@> ^P,O*U$_SCM5$_K)3NO C"TA&" ,)[*:'O"F_RWMH 
@8U E/M3M67SP#DUV:(G0:@CJ_1/XQ?(5@['\G*,O8>, 
@QT@.![7=\Y75]KB0S[KUC]//-\)W+[NWY\D.2>O[Q(0 
@'?N:)AB@_Y)(]_K=BQA(\.H? /8+ &$N^;4ET'2@7E4 
@A!"?4XNM,G,#5P1ZQF=6QA(+SGI/8X(< 8!:QA7Z0\X 
@^QY:'U8VR738@Z[P/<*77N"_K; VANZG:# .F5Y@ARP 
@7/2Z25XA;3!.0G3JRAGMY8'*E[5RH7AE4YHBN.(X84  
@I)$B<DVWF+)QBE"DPR!)6XN"*(F08ERPT8;-/I$0F$@ 
@CI@H_>6WYVQIU8=#0R%P;$+ 2'DY )YYQ69NLG*-D[@ 
@1NBCI&Z/!+ID4I4MRO,:MCF&@FQ++.<E;>U8/Z+EZE< 
@+'-&RH739?C*RFOS+M?'\[E@P42=XBLZ3K,4+!!O^#L 
@$UKJ^RI/P^W-E=" 8]"CO!G+W-_*9C%Q_*W[8WDNRS< 
@6ZLV:18IJ53]K1G;PR1^W;!6K7]^A/-;I$D1Y>5I>7, 
@J?+T^'<SP"T8*>D0) . >V#OTS=O,Z\8[\^C5!Z307< 
@@8-UUGB3>#!W0'Q!5S?(_#>5%]- N5[#V'4_CF&W538 
@,7QQ4 _<:Q+KA1O )^B*#T 7%9JH^U^:B@,4OA-60QX 
@VU3<O$"(&RX&:.B\LQO94JC5.<"F-R#@/,G9H5CK)(T 
@O_KV3 PE"0)-K$-%^SC:$X0H-YUTT+J$I-ROI/]6IW4 
@TATI1.E)D-_!DW*$4W@YQHO?X%S\71C*>4C0,ED=BV4 
@8A-%9$I>(S:>-/*$?F(J/ERZ;E!4"S'&U>4F-N#/M_X 
@3?82?%I8^>H<8K36&"\/K!32^J9=*)[L[#19J,I%WPX 
@WD>2NW_8W56HCT0XSI N30O=[;(#XIVNG9W=L&@%IO\ 
@Q5;>UVA_'_;*4J5;89GN^L*GHVXK!W];DOT,RDZ/21D 
@#]82MZ495TMJ63Z?6Q/[7X5F^X ESD_O8@+365;P/GT 
@[1;53<_;:6C^;1:%8<WDC/-67<?PB Q7QNKKTLWQ(&4 
@2\'0Y>/&G';*WBY+GYI9H"D(<<]8$O=WK^CYB(V%?]T 
@EG^;Y]TN/5 D\;V=#V'+.1Z[YL )4RKY$8,0.^JW7+H 
@01B=W'-$.]U^2.+DJ&#3ZIP$C*3OSA-3.3W\QL#*&*@ 
@,XK<\[(]-$!5NAV -Q (XE*2INEG0$RU'V"RZGI;%'0 
@<6-(5]T=.U"$I8#V6VT>(%O.W.P<XK2/<#KF0\32^Z\ 
@UW1EUF'G_QSWEW3"<C2T4#<NN#_APA&7GT.)A,@K,H8 
@S<UT#'T M'""J:YNMR9JX]H=J"387=5):5:6!F)XV\, 
@C4BS]%U4U'LA/#RQ@9#$JXD3UU7R1\EY4W=JOFD%E>  
@2_ZV;4FR@/D>\& HZA(S>,5OE'=@@AI::_^>T%]JXOP 
@12(T@V;G&A5VDI]V'K#7\$Z[TJPC?:IP?FJ(\<,VU?X 
@%5$]M#*62^I4I?#M %_\"B8+)]F""X1M74TP<CAP'9< 
@M*,DWI?0FO8S\CL;L:^[ZOA&MX8^U'B&>'RF*1OR,<X 
@9!*1PR+):"B$ *_?L/?."?^G7?GK344#I@9.(1'-TRT 
@KN?B<W--I02+Q5)N54^,X!=#5)U"8*ZMF9VUXYWS#U0 
@L'AQ@@9%Y0SX2KK/UKOS@0@J C!VW\?8AQ*G0F( 1O  
@RQ5$ (AX\'4!R7 [ T!_]MVJH7(;ME<H= &>[^:KEXL 
@,+K[<R4@!(WQ$1)BD4U#MO"Y%[*KOX/^#<<^'6X%(V( 
@?=S=OI%$,Y9]++(5X;K4&UGQA3+J*4P*5J8V;6ATFJ\ 
@KOJIY?']XD^53D5J9STWP<KBVWW;\%>B'KR($,])D!< 
@>(0+#H(..6AS_+SL'*MV<KIMK\ALJKMMX0WCDEHOM,@ 
@R2[49',3(>\'RD7LL^8.S*.ZB7>+SZ"ELS>B4>U"7^@ 
@U4ELRM/N8QN]3@"I[X:\V';Y!&HLWAL):E+_+;V.9AD 
@8+?SHK[NSFR^:C#9+H,_Q G0<Y6U\P/_GR3.75D1^B  
@"KM,Q*FQ,="P*>(/)G20[%YV!EMZ;]EGG);1*DVCB)D 
@!4>%9I7]@]*?+;CL%1;-BG/[GR01__&VP\A3G!/M.U, 
@%EK_R<S)TP@9OS#4;$9.-A-<KU05BDJJ&WS#_ATOL48 
@6U3E[! 0U_@YLK#GF,T9^W!@GHI-5-TS$S7T>[(ZB34 
@N<^)<8E3[.&C\E<T5+&H,CJ/DQ<DVV=V<8 JWL6.KC$ 
@0=G(WJ&G<8>7@-PO#2JKUS015<4II]>'NDKO6DQD>C4 
@? &0>PJ"=-*AMY&0Y+^@9_I$VP!!>8Q%\L!\4JW>S4X 
@X9ND;F<X2E %(*6DVW04W)C+QBP**47;=Z0II&%LG\, 
@_=RK^.E5V>:Z21K@']_@<;NBU>ZS(H<I>FP*^8ESP%L 
@JAF\ ^-OPJB2 ;/D#'3><RK:D=^XS?^62')R):8'J08 
@(3X8'+2.?$^R247,)"7?]/26RE\[5WY,5%J_,N]*6WD 
@O2VM EMV^T!RYX>EG/()=7Z1*EDD>SI\1?HB.>1D)?, 
@1P 6=VD/ LXR(/?']DW&L7[*ZBYT'/*7D\S&@%L6]XT 
@Z9'I1AE+Y]85]H99Y$;_1I;@7*O=[F!M&OQ'T^-7S\8 
@<?>IDFTFW_V;689,B+%U&J/Q'>_V<]KY(TN3;.^JK60 
@CDV+ZY9'Z6[!"]"A^*#XE='39Y][$QQ_-C 3CV*O,?< 
@VWX"12X%%#0:&1[QFK8 >4^TU;I2TIL5.C.J[(U[@O\ 
@SW8,[AAGFC0?$%*K$*^5_\A^""DA$:6-Q2Q8J5J30F8 
@2KM.'0A[++O)J @S?.:WI FP"[KU%YJR]-N>FLD+JUD 
@2BH$J'?XH;G]T:]Y5YTW%3DRY7?5<5=%Y1H:@_SK)_D 
@6S%^L)CQCR* ".0N NSYX9FQ71<2B:&4,0>TY<#$ ND 
@5CR&=9@B)>BP<!J[H34+OAM/("X5]>0D)=R9"TLOI,T 
@9#J8P%A+I7R'0SW.F!@<E9XOG!_:Z0O<W5ZIN4VPG 0 
@B_9NU(ZUT;GY#.'X,/43[N=%HZ[P_K"T%-V ]K"6("H 
@$9F>VW _&0NI_+S&9YCTL8/F^)>OM\H#6>.B!=-!D8L 
@;PVX]D#QTD7 +C:)@*\HW?'_V[KWRVV7(ITB@PE@O1\ 
@FSN1[,E0_ Z-D93+K(F&I^\U/HOF>]8+!0IIW)!H/9X 
@;ZB,1N*2)KL$B<)[G!?1;UQ&?.RU9%<@N%PB%): =0P 
@].!5>CUD[P,-6>'[F:KL"R%&1R"S!#8JM')RX;X-8KL 
@TCLI('HX0ZN6]M')LW?H$%CXY40KT8G@6K?+V7.U6@\ 
@6*-BB[6%@.XX%X<JTXS5X@PITX/-\O1O%C<-]?3?2=8 
@<@WIP:\(< 8CB:7TY\!G*%B7##T.R]+NJ#X2HPJ0:(\ 
@A Y'8' A7.I<.5N?& D%@71 ;4V(7QO68*IYN+7*K=4 
@FKMUK\&S33YH7*L6G-()6^@Q ?[@%:,S>5.FMF)7[SX 
@SZ\U7(=\S)6AIG>A.W"*C>*7E-AT+V1<-)*R+?'07<4 
@07P:PRG;7GTRUL=@R1^R7#R)9<_9E[\-)*?+%] C%6H 
@9O8;]>RZ>F3)MQSHM;-#6Y3R@17LQ<A.2QM_ P]$@^$ 
@[9WL%"4>5UO/*N4SC/EZ<3U=$G<XS5'"T,5:35^\_@0 
@GSIJJ2N.4 $L0ULC*UHU]?!56AH'6,:832%(+5V08ZD 
@C.W1.*^ F%%=OEP[.^845X3_6YKCIUN6#J-:O&** ZT 
@5L'XM]I)]"HD^Z#HN__ -BU1LWDG<#V\9\\ 3J6#O;P 
@<W0#V^^YW9=ZW0U@[/^$E9M)]>O G'=M3>^S3Y-?L#P 
@V)Y;%C9J1CS-:AQUF*)M:GZ:JUD3=[OM<Z1*MCD*,_$ 
@HM:KRGJ,4="PBT*H-!]@$E0?#[\)*-8*PN(+>(<WK$D 
@3US/OXF?LB#?A&?TFT!AX_!Q'-5UJ)0?RD5!=(QQG'( 
@ !!XP@&,+\@HC</]@MB)UL@-5^)UU8XUQ,MJL7=RUUX 
@F@L/EAA>]4N(8 W;OQ](3>+[Z]%983J;3U_X=LPXZT  
@BN0%KHYK;Y3#2T!(C9.P:3SMTSHDQ<2 6_PEN^JPA!L 
@2YQIYJK(=P8R%Y+18G6P=JUA_,4LPTOM0N;C:&(309H 
@5R$6>^FN<>=9C+_D./NVO)[D@F''A:;"H4H"5MFQ1MX 
@_VC;)9&5S]/Z2^1NM(YVY,?[0AG2G4::&(6G.8Y_SY4 
@9W.]J;:QI! F95P'X=P'$:\'Y8YB,.9SW3*X?I@)L4D 
@?AWLHC_9A_4<.NILBS/KZRO<AE5@'QU&Y0=[V=ZI[*, 
@1<8J@[K-1Q7 [#>^WLJ%3V2Y%[I* '3%Y3J$![\G",( 
@Q3/EO_>>L$-V+O!JU>$T%S[='5EHZB?+R"+OU%#J,,, 
@&C?N$NU1!YPS(OZ]<F'XM)YP:*0DHL2QCW8729BD+2< 
@T^Q3S6H+M\GE]K!%@/I>MSWB$A@MGG2^ 0KL6DVD&9T 
@]V,IU+ #"3]:GF;T*6I?T"ALDF@YG$MGN/\1Q)N=#I  
@!-Q S8$3T3L3SYFNS/"HO@PKY^",O:]44VV :SWSBHL 
@Z=F?W.S>F(.+#"KO8!P^-%G-JX.([3U\+;=E@UZ)LR8 
@S0?"_-EE.JDFL6)!V(]+%E-YII_;]<0EI5P J6H &"@ 
@<1?7_*C*6T\YOR'5;D!#U92<-S+C9E"W+]<'Y''SWK, 
@Z!;6^L$S]]Y #QP9N&1YQG%/HQ*,O\Q;A8U'#P5-=/\ 
@;#< Q&&C;["O4/NI8WK'<"VMI:L2,LC39_BWJ 3%9+$ 
@;/9>E$IF&-T9CDVBH6K2ZK[MIDG=[G[&V%MP>/VKE/T 
@,AG_Y-T+WX%HB-(M$%]6A<+O+U9;%^\F&-XZ)F%IC)( 
@II<1\9%,;N53QL<8DMIAH-,K$Q_G9UZ+=0DZ6V?1TJ8 
@UMAT>+EG<<G/9474'+"Y[&^F0:FD^HUE[D-KP?&8!3\ 
@,_@T&>%G1U1CM&D5E]Q>7/<WN!=L*M,^+:+5Q_"!8JD 
@9AQ!PO##I-4)%$5\9(AZ;#K5%-+/P*HUP>1Z SP,60\ 
@)O#JQ^VTN]]+O<U6>I_2T?VK0*)ETO6A5)S)D7CS-H  
@14:WAVUA$RV^RVY_KKL0S^SK<7@!Q.E%'7_NDRDD*<\ 
@P[_X=ML:_D/^R3QFZ)<_MHDK;DC0MO_^T;AUG]B/VM\ 
@PG_>[%13E0J21]HMB4"Y:A0UDM!H?=M,^,?5C',@H[8 
@(J9A1PZ.^<D93ZMMHIOEAV=83 *4>5R]3%)RVBGP_P@ 
@YCI085/1J:'GIL+ENL'?'E/E<=>:NID9N%_S'L$(Z8D 
@T,?",P2BPG@>7.I"STHW0B0$^=(.CP&5?E;>F]OG;%T 
@Y72%%7NA_W_4VX[:)O2*CT@C,U)C)R7*_+3FT'$%FI0 
@G?EGPT]BJ/2L8NSY_;X_L*@&1_7&]"64)8IUIXAL9IT 
@H/XC;)%)G1,L+]=LW'4TV48CTQR5S*59?[\-GK7K=,< 
@>LF_W;1%QKMXKKG8M[+PEE<VGN(DF'VYN@5KO8>>=<, 
@M32.]'&9!)W7/;.Q*$O_LB-.Q\VOQ2N'0(DSCNR3)-T 
@;!&A:?S)DX=%:PR1&XW*59K@A*X#G>7'9!C=SUF36/\ 
@$1CB4HT&G'$*,9&*<IR>"HLPXY0@WRI(&SEFAR=?9WT 
@CC:'0DQ8!MD.K!N;_79F-P( ^:(A?8Z F*"\C)][)H( 
@3W,"3^N6:HH\C67"ADA:3X;5Y7"XO>?UK '\1R)_\J4 
@;19%G>V?Q;7U4S20@9NMMEZ57;3NT?F(VCB/KGO]O]( 
@EL!>56<)>=ZGA3Q"IQ++;7U/+81LE]O)LP$FAJH#_<T 
@ LW$[]R7Q7D*[5_=>1@OOV1V4[<6CN!3;SVE[=N&W@D 
@@BTU#;X7EA'+%D)H%;KW0F[)'?X1DAD2:Q8.!:'IP T 
@'\%>RW8^] 7"=+)R>=JZ\^$2)@[(6_@&>) ,Q!>M,A\ 
@&:1M9QF/<=W& @M&F6OSUTBBE*OW]T ?8(L?<ERC!3L 
@@L;R).EP*#C>YJ)ZFGC0[<TZ='S+0)."XQ3S2A, R!  
@ZM]I[_!2)652MC-S/^QD9,@^-_:G9$PPB@6M?N N_ L 
@N$M4U6UT>?TAY[]-8;.ISY @/$*(.JF^KRZQNPVT-Q8 
@F2-I)41.J&WL@PTG3ZX4? 8"3X=C\7+$3UZ>F]$\(K4 
@DALO&&+(]@)"_]/_&I5\OWZH1C2]BF-UUTP&V.C%L%  
@^?0?1GJ2N/6U^KTTK+5 VB!XRH=1*CCZ\)>0L-&'B[$ 
@GB[FZEA\#3VS:UR_( #3U:,T'6-9O=-W6T"$Z(G)_+L 
@1%?O#EJ9P4LC?,7Q?W3 1D)/Y)^U-9'(&ES02TP=7#H 
@W\>YZ/* I/Y^3[3!:">_]>4ZK>K^,D4G/M!Q;5:.1=( 
@;@%CA:YA""=.2UK!R3;<3 RL-94GG4H0SA 7(O?0Z_4 
@>32); '>$02O[_>_^\$NY>'O0Y OI9<IC5LTZ-HA6%8 
@G88,6F%I<C=LE+!K4CQY+-#Z>/&+7J],>#\'L40I#C< 
@3S_P:L$R&L ?[F)AU^!16B.])1&9-QCP7F)<CTPD<AD 
@(.V63(P?MHJ.'$W45N0K62&PC%QT34VS:$_E.%O;B/D 
@PS/+/B?^& U]L#[N TPL&.V)A?-CF!5BFI+R6U1Q-S, 
@5T:2$K)&O7)S?"#"M/-R0*C_%[#S1R88GY_,)M9M5 $ 
@XJECG6JW"X]3F[PUMC0 \$15J%I?ML@X;^/09!?[Y*4 
@T)5)$T%[6PVH4 GT&"IG\M. DB5HK?E-S0V+4_TI]W8 
@:KE9O2('48< C00>9RMC>N4)=3/K&%R&"/EVB?Y%J5P 
@4_T6/%HHI:U)=O*4&AB+(@QO,@'+&-F:8>+TH=> ?&( 
@;SHK.C;2A[Z*/*>!;")Z'U30?WY]KS(*@M!A7=8(*F( 
@VNEI(@+Y]^:KJI3@>=U5,47UN>I@^>1_(B>'+=1DOL  
@5 E*AMSP//;T%4*_^51[8,5RK_QDK>%LQR=?([3$D2D 
@ ._4''*L\5W?]^4N32X;39C.W(,9L!=?F]'=PPX%R?( 
@ON<?$);LL!YK[< +[PH&CIS];G3(H+6%(X56)SBR3QD 
@>QT%):-.$(\,N+A"9X)/03-:@^:2.$8V\J;KFBVA][T 
@L D(\<97)=(#B]:)O3#&[#8>)?F% 4?U7FQ#5OAU* @ 
@N1#AJEBTJS+F(FKB.Z%*8[Q.FZ[7'HN)V($4MW<QKP, 
@.KF\H3,FQ((:E7AJC85>$T6I3E,W2QGO="F\&AV8SA@ 
@/$ZN+E/0]+/GQ&,4@ 3G$$<^(H6[D#@/R;\)@1H%-*\ 
@#YNH(@F43)JRS4IGN= 3.KC'H4(O-2OE7\?5S&ZG*3$ 
@'.U9*KTL'"%[^".*CTMDVSS<MHE#4*) 5;CRADT*'Y\ 
@&E(2$8"KRWNS)9L7_B4!D3YE^;  "KVQ3Q43CXG=!!, 
@2K#=>.$KC#0 "(,T<@17!<(>\Z+D ..C>"]@9,:XZ0, 
@K9;KR$>GGM:'.\AN<JU%]:S<LFX1]T*S+@&S\27[I7D 
@OV.V,I\X2BHFHA-=U)-C<[2RL2P*1G0,QJWD,P4DX68 
@U]S!1:%UK?9VBPC6-F,D;-QZ%7@18]IC$X,9EW/D(UL 
@QER1*#,-&68%\U "'S:J[5CA:FE.NM&NSZ^[<I[^/F4 
@+">)I-U(/4OL>2Z EI'$1;I%3$NZU^&-\$YG5RX^-BL 
@D%AWB/6&6@*?(?%=40Y8Q@FW]^F&>V=@H?_E9UB$T\X 
@-?+V(*FAKP.G/#F@;*'H?;SSI%[5)Z3>H)1*?%V!1DX 
@\*&VZ_7<,J<JSL"D=!L,@]WV&?V]3P$:/# $68HK5>P 
@CEBNY266:!+?MOVTVEJB4$($LOZ85<$3I[VM,M!-^^4 
@Y*^(^9>8'?NV(^]WY1I7H<\3RXDQ27M+S[SDM[7QART 
@7Z[[2;[X[OD"TVT$7$DFW;M>%25)L-]!_W9I<Y<Y3>X 
@:")G(%.L%=8.ZF1R](@/V@,1DP3_826\3N1#S@3TK$T 
@[,G5=,N(N=\*-^> +[ Z8*/)O;B8[>]UH6'18HB.[6L 
@CA8:IN"+,U\M[I95+$VKF>Q*;+MIXCVVX$?XXN_ZA_X 
@D+X7]M3.[NSDS)%FGZ"51F([FXY>V3N'9.3"\D.WD9X 
@X7_QQPM2?RI3F(]"2EVD<)GNF-6\M-P2(-&K/RH41\, 
@\!FI:).-L$ .+L4]NF$V(-Z3Z@P318 A-&-E8U1:).8 
@B?;+,>&)/;]+H962[ITKD/,J[\EJQ9@Q:2MY#0+_<*0 
@RL7(B(SE(4L*^W!L7@<QFC0WG< 5ES)O:YOH7S#*3A, 
@:V) >@EJ8;1&(*AH6=\J!1$$$HS@8W.0E7O*U1PSVDP 
@TX7B<U%>+[U)9)<:)^<EL=C8)RH6VMW=U_;K=2Z<]14 
@-$X,K0:V,&O7YWGS1!V#$Y9[>8ZE[;>0GU@<@B3$]\\ 
@[X2@@S^3*@?A19UP(\,);DJ33(>JI QE9OJUN"W/.;0 
@@&%B [1T&&B#/]-6/M8'/1DXCI6-FL_YZ[[Z.KUKW>( 
@"UFN;O-M?^PC$$$L?#LZ5!C#1(]43:"M"80&'F3P;7< 
@";8>+(*F<)Z8P974<_.D4-2?EN0',#6LH6OL<I=6?<X 
@Q5T).H_U9$"DA0L1.*W&*70[0=C$&FTA 0%*$JB85H@ 
@/8SE#I0"+#J@KUUA!\@*/#G+ +C\(+.G=D(O&>LDOTX 
@"Q?C'D+"BDV]!TB<4A]]M;2U=RVF*7S<]"I=[>L/?>\ 
@9A< _NPZ5:>%@6E3#!7YG).PF<[1!%2SC$"ACN\HC:( 
@]]5(&]MAD$:F\&;7V^&VB?B0K<2+PS22F%"F"8/,YG< 
@@Y8-%I939ML0N,B=MP\GN-JL5IGD<DRG(#JQ.G5/Q0, 
@!,_BHOZQBJ2*\\@A<GF=,"\U<VXE#)[).?UJJN!NL=  
@-.SH;"B:LOKMVTVNP\\R;MMFW^"#^80OY,D/#+916,\ 
@T/,&5 B_+0,EKL-DBY#?KOT*Y384/J'TU285-Z%([^H 
@X%=#BQTS89</I]#,<Q5N^#X1:=]G(Z$Z'&REY">U*4  
@=YU#G^%]5/O&<'%W>T:6_P^U#X_=0PYS2F2CMR05%&, 
@OC7[YMTK@#X11&6KR&)*^L> /GS"59Y50#/C%S+<71D 
@*!4%-E41@6B%/)J:2\P/DQB3DQF31$S.Z--3]:+L*PX 
@R8W[WPJ!UJ?S&[%$A$T@S*C/J?F^6@7ZEI<M=$2E8Z8 
@=>CBK11DG& ]MASKTLD"X*O>2C$;G>:69VG),AZ]D'X 
@K,5<G</2J]5P^+PE QE8<./,P@U+B0AF6'[$M7)<NQL 
@VVG1Q63/YIZ$5Y\!R=26@DI->;9^:4;S2^?U1%9F#B4 
@X&RF8I#].XSX9&99^][HP9.53"Q!I>+$@_3H#ZJ.A&\ 
@7ZT.>K*#]DK(E\@I=C4,W(NA[)+QZQ[!^('0QD%IN3@ 
@-BK#,G8_6Z\A46=TC8N,GX. _<ZC,SZ<3KWPM9ZC8B$ 
@!GUEI/;K/.3YU,0.WH!DK>C7G,'6C'JKU'F@EMNE^P$ 
@A;$K+/5?3)!HCN!8N(5<:_I,6IZA'#<C)$R/'UUK:K@ 
@"@ 64"SZ9.8&"].#$[V\T$7D]80@Z11+M\,786#8]J, 
@MIU[E2[>"F1-Y^X'SU_M1=2#D"[**D/C>,41A'UQ6U4 
@1%[7(K*H&[<"9.$#9?^AE\DTI-<K+WE7=/K#%\(G'Y0 
@E%98<<RWAPD^=\Y"($5#VJGTLT!BZCW:=3W?=G57S%\ 
@(W*S/B.MB)>>P'<4:YY;]VRN]#R_ '[UCOX'-40T]7X 
@8ILLE:/5T$2EYL(0\&M!RU(7N#L3Z(845O9LEWN;L], 
@;Z0$WN]'FS&0^3N9F#_8+^>7=3$F#JI_)2H=8FM!F)X 
@95>%V[\-D[&]?X@1X.GH >[$+C03=GFT&!V544I\5G, 
@&B=?1YY4(7M3$@C?)/#Y8R*#KU'49>#84MN(>8+W\4H 
@?N[V$&(H>-L;7UGE [LH,M-PV57$:@RP2NB3O&.M?2L 
@<*S?S3]C>HO+Q,FGZ:^IV#[$VXYBY)IX5IKT&R86.3D 
@HYC7^PZ4THF 8C%(+21R#>.6&6YN,4F@OHF1]P%'#@4 
@0VE_; ^Y,+1XYI2"25$#BJX:&'?+I6$Y?O=AMO)EL=  
@,LXV[Y6F+EE'0\]?30*S+VSQ[6KR(\^W@SL! &)C#;, 
@:TU<4'\:YG\205CSS_J"L8\W!*!\@+*]'<Z"X'F3280 
@\//@#&-T@I^!#R/::YI?63&)7KLL0G#E"3'&ON.Z?(X 
@;[Y--6?FX6[ TPQGHNK!>W6*1,"S /C%CN5?)8YM@)$ 
@>4ID%'A \"!H72C9,%1-K(.W;C.'$]=1I&INPDSSMTL 
@J4B<)3\6<R6(8-\29_+"$%">FGIK6-3IJ%TWY)37/[@ 
@<%T@/[7J'@1P4?$T5Q+#3[<?Z20F%-+UO@H^-5%QU38 
@T)RV\W"6Y@Y>-TO:31X'8[E&B@[O&+4C%+Q3L_C^N^@ 
@ /T:ONIDX6],W0_8Z<Q^R_E\>R]>"X]0P@O="2 NA)X 
@<DB@[NAUM838&2P\HGQ<[<Z0LF#=R*0HD*Z7_#&"S+8 
@!A]HNVFUUQI0&9X80%H1-)J@5C<D<NW:E76%;:@!?74 
@_F=V#+EMX)'X9JHXK[,J.AT8>/#H-?*W=B 10M;11(T 
@/:7>:E74\H]_K!Q(_[@%&"/<.W_Z)E]Q%(?U,#WOK(L 
@B5@O$^>N3&.K(,GT?,%3C)#=Y38ARO1U<3@02G_IW%< 
@)H3XV;&UP__&8/U6E*KN.7;J\!FFU[P'.J6L1\$?JQ8 
@5XCU*Q-EFSMWT !I6!SX_F\*MNKT8F P=Z/<)%8T67@ 
@/ZRM;HCHV>%WH )H<"LI%$U%/5+76K"P-J#()9$4@J< 
@/3%V1]P.JK\NG'J*T7]&@;Z^8#<B^R(:DN52!K-(@F( 
@$B_$2F">6Y4_23_+W3/V%LPP:ETP1,DY. G@MU?\P$X 
@7)SX=HKD;_>$,Z*%92,VHIWQLQ#SDH#U9@D2\7NZ!)4 
@]^OE?S'53Y?P[H#L:DW<^V V:!* #Z)=%"BUCH2>VY0 
@^FD'0@XW]4^Q=_E(/HYQD(/7AB(6\3+3+B^X7CVS45( 
@6_&OW$#_ K40N!"$_W7B*8,(T?,KYX393INXT$3T\8H 
@^&BA[_0QS$XV^VA/=GA*-4NX^,,,,!\9R,A;_[X[CP0 
@,<W4(Z<;\#>O_?#W5G>D>TJHH5T?WUTIME_%;> 1EC, 
@B@@Q_BU9^NU$YKJ)F$^7=5#BLF;:\;M[Z<[/%I&S,1$ 
@XD5)H[-N;:# E_GSB"2?D",=C*,[ORN.S(DWG>?M5-L 
@?E<L\W3%@;^4^8T9KB<&<-@Y"@OL=>0EA.37-_,PO&( 
@_6S:E"D 7A8\-B,S"_%7794JU"@142R-BV32[_VO=N\ 
@R6H3P\1H9;(H'BXC5LT475_3;SJ#V.$WF0O\'!/X+"D 
@(@B"W5*S191*SF2T@%V<50U1#*K/KIB(5U #&'/ZBRH 
@MA9M#JJL4^'^%V$6JN0NERCS%YI>AW(BGO[3?X$>-EL 
@99M#8'Y/H7P!I!!DQ:\N9--\9&,K<5^N.WJ\A3/HU!H 
@2F:G+XHBQE?EFF,O@#,U#RG\\G&^[_F(, NRM;'#<#  
@R3JA*ODO*MC-\&7\+#SY6K]8F55_-PV7A8<TL/W06J< 
@6F;1'3$QC2U'HV2ZVZ%A2\GQ"Z$#]0C^L85M!/2XTN\ 
@C5,CR+9#W.%H6Q5Z;Z M>W+$^&JI.7F8<#REL[!8Q=T 
@.H*_EN0]]N4+^?_H Y!>!6\Z\5,J8:*8!=7L]C@DX;8 
@WFI9SZ<SVRV-9*R46G+[]VXA_ADJH!WIQXF+>+P4E?D 
@-YJ"O$K*B!UKE@PEA>OQ0Z[I.? 0\@F&DCGF'IP,S-P 
@Z/O3#M)3^KL#/H/.4^2_TYL0AMSU\0_M1TK/% 6Q05  
@G.,]]4//_:#UV9K.%1PF.U/OH]8]4IMI7/M%@WB> 7\ 
@>R-#\?)Y:[UY<*?:N:$6A2=9",=/!]#V.*SD/ ,BZ.  
@AQ[^0UWH"4;M8"CU"\@'E0E4HG6[OD-Q/>**%5_S%*$ 
@QB@\U\K%PB4H5+,!\9A/"H$[5#34%P,Y79!^E?8M,$L 
@JZP/V*"J_TNC5?SB]^I8A"A#\V/_SJE3 FD<1K)S6=L 
@Q(3.77H$KP'B=6"3G86_;"L"6;N(R&YPKJIK=ZV%,=( 
@;5)YT=_A.#VR4 8L*T11Q[T VC'.]Z7_])E= Q!+"9@ 
@KCGBVM#/J\!M/\M^,@MD9'B+5T;P@0F37'Q1W.2]A', 
@ 4%Z> -'9Y:":2;<JR6^FQ]LN%A&K?]1(ECGF7!?YDT 
@QB=Z%X2*#)NVEO)TBL?IE[^C>*.^N_+T;E\HGU%_!Z  
@H $A"3<LU"'G[I#8B^']']FQ,VQ=%3!0=\3U%<J*.G8 
@P7/S^$'@B\ HR'JDCDIZ8)LB9+?=.EX74UW808XQUFH 
@]V>/P5",9/-DJ98# 2T[V]XCIZIJ(>Y(H0ADO(LSCE4 
@L7T(I)1,$^#X^)G+ E;AU$\A=.;7?\UD!C4N&$F\#=( 
@VG0"?@;Q@Y0#*-#>N*:DSCC]I-:AV:,*32'40*94M\\ 
@ .)<.&S]IV7OA=XP'5VE_>TITOZ2Y*S0H,\0J&=#C=\ 
@;[;,;L;Z6J-8=%O.7(IO9R1&_'8[O>HN [>)PS\SXET 
@61M^HF) X]CKXY4MCV[Z\EO[(8LN@Z]])^2CWYD%#IT 
@V 'OZ-&6IT:MT"*0;\$71G6!XOR3E,7-M4D-9_XC+I8 
@(7:W->*R;S_":B4KYZ1H&%M&)#JYB@77W,#P8*MM*88 
@D%VH"O_G]YCD9-I=0,@73CY)7FA?6U1+I\F=96Y$%SX 
@<68K\]4]0"___5RHQ8M6Z;6'@^B_NC94-B?S4O'1$O$ 
@K<\%(:1)FF/;<'_=BRZ3-GGLY@,*HUM+5P15QE%6P7P 
@ $V#(:^/@"K3+SC;M_I+ _%6S$$;K1XUBBK+;).><,D 
@PO1@]39F=2\H[TJVFX>U\KQ18FV9V[/D6G0%S>3T9W@ 
@)C(E302S'4\>,,QS16[<( <2_BEV>I*6FJW_/1YJ/F\ 
@#D;C@3W&$Z<-YF4]T5@&G'J;ZTQ":FA.!$C_#W@V8'L 
@[H;EYJ@4J21>8;U& CTEG0#0PDPIXX?AYI4)C7NC:@\ 
@7LH**+DZB!#=U*\" @LN00:8J C4HQDT_4A]:S,-%U( 
@IF[X\2OE^&XNM4HLDZL4Q(7:'$>J.+6SSM#2%H:F'6H 
@[OY'7MN7M^-N@M2>R$L"HQ2VYK>3W"7KR3O':" EN98 
@WZR:?ZQ1@Y]>.(22A^=7BY""W=-TG=YA/^DV.AZC>6L 
@4J)S_!OP&&0&3<W9?']&:,?UQ38:LF4Y22T(.,)%(T\ 
@IV5A0692WJ%$C#2J+,E727$GN+$P, :IT#>!F ,!QV0 
@BEM\G)H[7#Z"?KP#7J!Z=+;F\TR*FGX83=@.QM](ZV  
@R:KLVQS! 5,5K&F_PH*1!698G%*VE:%REAU^<D ;<9D 
@V[% "B!<ZN[$] *!S.C41O;90M#384\ZP]V.<&=1K$X 
@P(Y*RA>?Q(*70XXC.LP3"M)3-#*5<*GE=;(L0Q58/_T 
@^E1O%>>T&GC^)0JVR9U1-^N4NM"8*!9)J8ITJLMR+.X 
@H'YHN(A&;<=A>^]X<Y5>OH4[DD^1ZHN(KX;H\3SK*B0 
@(BNH3^[I13Z[ZQ14]X]W>N(BN<Z7&9PD:D89AE*%9F4 
@?&6<O[$]%H;%RF]S!PW]"]S5.<@>)\S.Y8I;OK8QCW, 
@& 1![=>=SWC.H$ L(EF-N2T*(2/EN[2W@"9$=1^$A20 
@T-Z>Y?FC))M$4VJ#&%N_A!G'^34-,F#^]AV:F=FD!8H 
@!DN2&31,.0Z3FJC==*KL1+ZO/16)!V)C[N]'$(X971T 
@&O <94IZ9W2)SSP(79K2G'ZE0HX5LY+8,ZWT"PV53Y$ 
@KKSK5]CYN'ZQT<^2Y0+4-)45U>UD2J#_-T8VS*O<!D\ 
@\@+(ML9ZW&L!:#=TM2/Z:L:M0F\*>!"@V<TM53$"#1, 
@C"\P!L76"$^EE*62,8FGS!PRGU5TSZ* ]I>PV'WM/4X 
@=[O@HHN^OI\D&Z+6:U#ACZ;DPEA;I?:!%?#+"G&^<[, 
@2L77,FW=+:5G.,:KS&6D!?X_F62 #V/7C"0!HDN3Q-X 
@[RBPC^(SE!0;5;>OH<GP+Z>G)X-$4Z88H0A2Q? @Y-X 
@:_),42KV5^(0+8M7Y@S90N_=+AE1!UA7*X7\'V']/S\ 
@[=S;!5>LGZ=1H/MFYE>W(]ZW725%H[8Z C5Y@>V\$;4 
@WQXLC27-D?CEGV[.J5-].#QO1MI9-2 :R<CUWFSCRY$ 
@:3O)EWT9,O_P$A>U8T^VL\,X9L*(3_/-/'=-4+1JOB( 
@.I%3RO2:*XJ[U/@ZJM^1R2;'G%%(;^CL8 _40 Q$G&  
@EBZE4D=3!3#8N7"LJ.TIYI0_(MHP,)#7TV [WJ2<.IH 
@^DCU'H^-$GADBDN<Z:$>;Q#2D@^F'"S4D2D-SL)V_D$ 
@C@U;]<YOB3.*H<@= ?Q@-+TE3I$['WNJ4,^QB &.F&P 
@(EY"EOY_ /QSSQ.9L86YKU#P).&_ZTY'SJTJT20=W?H 
@4S8S_J_'KCWK>)_:N#1ZE!\ I9\L')VE8N!^$KK;"]  
@RI/]L]G#SA3\L-JDL#WG\O95VA\Q8P<+1QI(2S^^MCD 
@V$$6 B8 TBKAWP)J8]0TV F,<W$CP8@K.@HLU$IR6U$ 
@Z0L][9@LQ;7@!\^>P8:3KJ]N 6T;2_$5I0$5U-)7?D4 
@'2JF?#VSH&]==OHO7APLH)<B"**H.@KJI29R?$)2M)P 
@"(;[]T#X[LOL@T+AL2 /BB.UHG;3K9L$I/K83W'XY1  
@_&AT)=5_.OOU:"8(2=&R\:S5YU@N[W@5.;=DN @:EE4 
@%B/*W% ':'5^IW<S,1?U0AR?:A"'(XU/LB_S6A" PR, 
@ADZSMB$D*O:]:J-1,*#>3<D[[248=.<X[*\@,FN/4#( 
@<;T6@Q05PK]:_+C]MR3']):&.<L'RS<0<X>LK)&J4*H 
@%Y!Q:K'DHT'K0NPK,&Y!H3C6!)E2U"R8@$0$45NN-B( 
@05H/UHRU9 YM> ]= 1&IY0)A3*&08O+#Q(=OP0;CZ&0 
@A>E[00T-SY9AM-LE@U_ZK:4$B,Z1R+?HVG'Y=7%#2V\ 
@I\]^ZZBO &@#NN7A]U;G7:]CO55*:Z;$5J-4B6)C^?$ 
@6*^JJ^"Y0/K@N,X[K&\'/&0TCIE@**[?:2QM"?'ZE4\ 
@>=4J!.+B_RTQ86V\B)QYCMF'T-A&HIE:[D=O"/ZF*Q0 
@M0S>;^QMP$EHU#5<J_(2R9B4FI;NACD^PY\S3&)J[3X 
@Z9.C;)T-FWMYK]OF/590SPQX_!_5[]ON3>L,"?G!!4P 
@])6FO3#R5=*K,=1CQ7Z'),W:G$QJ][(!<=]6,D,.T[0 
@.Z<D_RR;I7$['&.WGD\C5%', .?4M*!A;G&\U_6C; D 
@<N"P_@RRPO82$(%/60=?QJ Y^C-2 YWFKW5DW.:A R4 
@%6Q^\5*2PNS/9BHH?QB.K&QMT'NXO8L]4-*F?P\J2&\ 
@"N<G;9IU:MK_T8UG0$QRVZ*/X('9Z6O]U9+6_!_F\'@ 
@ JRFBRAP^YW9"28L<N3M5 *NDJFV$:&'[(9DQKFP._$ 
@5"8@F(U'H<QXCG6$('DJ;I_SL;\H;,H^&P#1TJ; OI$ 
@VH_1WIM#](E/U*-E]J.ZKG:DF"?9-;]:?L7(%F+UM>@ 
@Y]@(,G7TF:0-I_8FQN/0R:8NN!SP%0U*4Y9LEG\$-K$ 
@D1)L>G,C4DKEEQ:'F9P\\8;L@+?X&$@C7J3=[Z\6 5D 
@($UD&!)J\/]KYEP=?GX_B7S?8^YDIL92^ D75N_Y5L, 
@2L#TC8[=X%PPN!V9G67;K8)+9"(^2L0W@%H.D]<JGL, 
@>,4Y]VI,\[Z#4L8KJ=#J]IH9M.D.%!PA,)!$?=].^70 
@R-U(.K,[FOJ]J0?P'WK=/K_<BE?O8I^74:T//DS$J,, 
@6XBZB$DO$8TI*RBD:9:DH''?YDG7M40F&M/ZO8RQ!GD 
@_F**32@T)'C[,)2&NWCN2J0X8H+=1!IL#4'7_)F1I\X 
@=N741AURXEIL^>1$V-;O=&'<^/($Z<]86)Z;?PRNX10 
@L7L(@?80*9HK-3JY@[4S$N^FQLM-8["Z#W^HI;&WTQ$ 
@G[.R*C(*OBOBSF/F1_NIQ8?R']%B-87#5/:]..#A5D( 
@OOW2N[DU!^@$M+*[;W5G_ 2K"\^'O9-Z1CVAQS)1  P 
@+/V7SL*R&IE)R@>Z^;[:$%S=$=/-I,16LN6M(O3>^@  
@W/:J>08*:C@*2[)9Q#M+FOE:96>4U+_A*86>W%RI&6@ 
@'8<:"-K%P>Q#@^IG9M\!UFGYM':H[5;G1'A0$6/SDG$ 
@VNA7'1*DHG.6592S$DIR^S."(91'$],G7'SEP2#9A,  
@/S8/6A9)_S^[8'7JW/@?]E,D73^(.:8^0%1)3%-.X]0 
@4?2[#PX,@YPP&)0&%JM=8%[U2O8?<J'.$22N%@U&A)\ 
@,&^W\Z;P\4_.KE'& *I/2&,AJ5394T$VB\B25EP.66T 
@3&_6AI1CE\V^ 7X[IQ4ZL@OJI7BF\@S3]WBY7L[;K7D 
@^1!$PY&Z+1P>0LLAYC%OF<6Z@'1/ V'MIST7COB,S@  
@;36'):2(OMU-&\<8[_JNE!2;4 J'2Q7U_61A:1^^%(P 
@,Q!>?8>08-T@L/B;*IDC+Y5(1#!VM!4.%.EDK<LG]+$ 
@OY70&^WE+EL!%X536[41W(GTJQC)5 ,A+M2Q@AE'P"T 
@CTX8"+:/5*E_5K;WJF51*?_19-X=U\0.?#V)2(@-6)0 
@OE.(#1_K+Q**\L33[]J3%/+RB=5/$)0QD$_RW<;2.%T 
@KVE^4I'*0JBP"Y?%NGL9/:)H67VOKG&?Z92UW3+@=XP 
@&UN-E06,Y2/Q#/=_??^3E,(@-]3Z4.6LI[1PC?B0\]0 
@CQ /; LP?3,LHC WCYOB[4#.ZDC\FV;"D#UW(]$N >  
@]%PZ81_N N0O<M-I#&P/'7V<QJ2YQFR#B*!K@U9_DX, 
@85'SY?Y/R.G [@,[83,RJ*_0#\9'9AO-4V+;(BXD&WL 
@)ME--19^UB!.<63 "ZKNJY:"XZLO$F_T[Y$0DY+!9<T 
@FDE"C*\98_K _>2.'D?:?3H!_*QD/5]%Z6L![J>3\:8 
@(>=T=,/SA4>6["WJ_/$>6.<Z3+,4D$D'@KODUG]+2^< 
@N-)XO>]T%C&4.R+I\+K6)W6NB2"UVK6?_$N1K+P2BR4 
@(YRHPCD(4+PUU(_"O):5S3S.Z9Q@'G[VU]0ZJ*"AT-( 
@>$C6Y8!5'6H;"TLD"E[Q&$GI'0,#/*B55*?$I$*HM3D 
@[X=]L N/X!41O[$#3W"\'\4BISQS8OBJ-R639.7!LD$ 
@!X,/P8<MFJL(%NHNXP_Z-T6TS F9?::^\#O.$&2:]U4 
@/TLO%[ENY"3"IE$M;Q.IMD#R].9R!K!@C7#P!H0,RM4 
@QSXG#!$HWL,751@RSC\3H39*!00*,IL[. &2;^1- %< 
@JO]<:C#N#QEPO-P ]M3 J*7/>93,R7<&(&9%>P#SJP( 
@T+/_E0_4.<I#D/5G 4_02%Y4U[WB[J<I!68K0P&$&P( 
@D$CC="]-^B:&GQ56_1LC'<B2+ %Q-]5EK32N0;5EO0, 
@!*"$VVU@;(^N*QJ8*(,)./QH20P?\B@$ ?^NI;WASXP 
@J^:!_&4JW2V&FY[*E,9IK?H-8'\I@TYN@)\=4D$-"C@ 
@M.Y6S$8Z9GQP]?\P\&1M5B$4L:T#UBMM \ES.OP*ZZ( 
@;U+_8?PBW4Y*OGO(M]X4?PN5K$PM-*C[N0[(\BFDRZ, 
@"JG A;I#Z"DNPUI,-B#@9NVT\G"X#M<>#/;F:!R%*V8 
@4 B+O@8T!$+NIQVZ8<+CO(FR)1*1WN>::CDGBCSN%%$ 
@$0RG*@8[TKAE3/!*+6[40]:BD-U@G6)PG_VG"\2WROX 
@N+.AH;1&WTB_\ 1_? LJ&80$ &]]VXDQ,70X/[=%I.\ 
@2"B[SD)V;RG^(^:\UG1'(!EI<%^N]4]^RXV'$Y1)'OD 
@5Z3FRF<J[),!*CS4*M5!$-E8#7); 0+ZF4Q,SQ6S_"X 
@/[$"&\XI/)>Y?H?K_XE$6(ZO V+\&]I'L!*<AT(*];D 
@JP<-BJN+)RTHC;.#GXN,(20)02.P>_2T)SYPAQYRS1, 
@SPTMW")"[=</#@:M/8"?5R7$*T)?X<X:3:U)A%-%->L 
@X"I0KW4TC2OYXJBXB)X^(9>,,OH2VHABDJ\>.!N?7MX 
@BY3%XZBI=>@VP+&#6!Y*18/>?"6M(7T!3QMVW*H0M94 
@+(%]!EFQ;M1R@280'8TN:HH@33761_X!6KY+Z:_HI%X 
@S@-/G*P\GBH3P>/FZ^V,+7DP,^6%FIBT2 &R$6WSD.( 
@'7IN+/G,Y0NH<(:^!5E*"[.7"'GJY^WMG_UG06^N0)L 
@HV)N%>U!JUL=D!<*0"%2#X3>D2Y+]69M3.:-9N.V93@ 
@MHH/8KF79E&&Z[E[3E?X0$$-\7\B\F F-K:.%*8E"TD 
@#@%W^/;B5(=O]#NJE&"N-]QF-IH,ZIGKQG)Y@ON^1'H 
@8OX'1*R1NT5_6,Z D6/2.V2)4]#(/Y11A=09G<\8^9D 
@,7,7.@?=DAK?,Z1/A_*3)1I"V@1LKS#=-:>?CT?R$74 
@A.G$OWK\I^E!$S_<AC ,V4F'F. LB*/[.S-E(BACY+P 
@&//V._NL:#,%(]M72@/77S]RQ*]OOOQGU 86&;H-_AT 
@FI[NE<G5I&(41[^WAE@P:M 296B!&ZLK >HXHM,S!J$ 
@D>D!NJ1K[#Q\Q<*I_M1^( Q#HO->BZJ7HP?1Y8H8[O0 
04^+7C!.-!A((L.N*RI EA@  
0=FJS&6WZ4T-4G;&=7+:!E0  
`pragma protect end_protected
