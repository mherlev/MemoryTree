// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:52 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
EL5jxoqC3haChc4B17lyTQbwEcLl4aq76oHE+imdklTGS49Pz6sYeAmNlRAJ5fe8
4jMmCoc4YL5uDE1gqyRXbU5BLwpXwBTt1iObDHdP8X+uejh1oYNmKUDdyH1KsUS5
8ez1apimRG39aZlR6DdqkBy9Zha5aKVcLDkUTwYuTUM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3312)
IBaZbJsRB0qqKDfDHSt6JLnqO41tmeeDq+av7nTBUYYfyTd3Qs2ic2BzEnCMSlEx
0kSdaxyy8z6GP2VJFJh7dGJfwzPJEkmJzPntLTQPheJHHj1LF/Rz6deTLZBNUP+C
mkg8v+7Ujy27OYmgCzPWQhu/QgD6jNWpMJDWBSu4HevyOOWuQ1dS+KlvsnCcnk5l
DiXq1D3toipHcDCBQ4LiVOmcYO4qv8NhQhNfRWVULYB/NpZm3KymLhx3MjNwPk+1
+jcgPwam/Emxz05VvXlxmT6XoxrYIDHyTivzpSVFOdAcHJtITCzdjDPZV24CagaD
VSlebGA2DM7gZfkpZ1thA6DjVJp4MVAWkqKUOGavx2eIq8VB9tH2SluZespklEYa
H1bNUHbJd+KseufCZc0ASdZIJiBq4g9/QOe4IGjmuZdrHyMvntfIb2jScXgJai0A
ECE3IDHsEPKBGA3QswxTa/Ypq5wLZj3kOwajitPp7c5j1NGZOTMnu4qU7iz/dhuA
aRg4XkWBKzyddy/maYA3gaOC2XXpALOekgLna39vTsI9bI09mCWYna7WhMuO9c4r
PECJE2yhpowcwNy/vuzbq9pSuNCpXqpKMiU91Oj54okmUuxIRfqWNnyC0ySXH0up
ZGEDog0zoEfOg02LzbV+2bpYR08RqwzaBxLFZfM43KVnIOJnnrhgd6ckmSJMvcSf
40vrsjpRjd+Xx0BXa/NchVbF490nkb2GLXNt3b/pwuh3QhQ5yYWQXjQYGNMWYplL
2Hh4WbgcCopnNSLvt62yOlnR8GEe4WBzRaLXai07SqxHVGFbs5aZPf8gheoq+DC8
q0QxAnkeANj0qhBwrjvWNfLPJw07PgJTsbTM0XyN1NEtS9aozncthNYfOSFhvUOX
x8nNTKLV+E1tLY47prYt2hXg3ru7O0ok2ReMTYi3mrnYAWZxI+cUZesx0mGkSTKH
srOfhRZUf79PtVYWHFiTQA/fGSo8coIPEWoTGIfjJNPecCDcNavsq/GCpv3jb/eL
QxbZqsfe9mIP+ompY4/tBstp03NfmehClpKpKXADIv3FrbnCmLWTLrLFu+JBibFl
odQC8LOXg8XpFj4FZMfnxIC3xRn9CIdCK6KQZfjXxySXf+qi2y3ripjajxec4KXA
ZftDhrbfQkLAQipv/t/Og6b6/cCZvxEiv8SEy6HcIs20XieyWjg5fGl1cbjCHnle
/XAjfac2xGUsBgxMqvqwkIxdYp8oWKEXtQfbGtNpWDSYEXbB4liJfAS/NjILLcMJ
rl1AKBuSxQQ++ISg9XquViXXo3CJLOSML2EXWEIFIW1yPnGnrM5G+AxT/KQUGx1r
60TkFqUrv8pPG7Bk7sWRAdVx9PN7I8q0OKfHWQF/FUNfjKGSI8eEo+JJzAKyvts2
tA+YfTmsHsRMexchHpGbHmRCeqlp+NWAZn/L7CelsnlAZPy8CarcJL+VcCq2D8d5
jpVnHal0vI5wAzc+x4DKfknULi25zQ4aOBWqbUQsCxRCgrT73vZFHvWmALecpKDi
Y+AjiHUPcvFl3vCLLQ8y0IxNKjtVf7H02exhLVJvkgDp4mgO2w0k0EcA1syqK5SM
RE4qrLN8EXSlzi8/WW3jeeY/ju5Pj3JZJycpgoze5vIQPJvhgKENarqMc+2YTL3r
TaTCoYgDTkwDMYacDEuxrmhIOrexZkDr8n7Nf7rnBMa6noncdC5NmbDkCPhMMiOt
ZP2ff2HHE4/i//OVneDRGUq6ZCbPOGDwCEuxxidOQSyw4tOnxc9O9MIX1thOv0Oe
tCXazWQHLfH7s0pNLX0ua63ERIgRetWP04hGtOaqb5AZLW16ZC9LaxHoG4yEKpSm
QHURFZLMk/u1BYfi4QrKtVqTRup3IhsSXDrmMhSa/TsUpHtAOLOKAO9MHyFIw+aX
6F5oxacXHfwPozA1N9C4oIvbDlzkePnVLMJp6R3Umvn7ZetqUH3pcLfubygGLGGP
OYoA6IXFr3Y4UCIfNsnEaezWogwmI4CQQYkgL9akhwGjKZJBL9fHHtptPjzr7/81
Ld+OWhmKu58E7aTyPf3OA6gXhrsy2GWgVK5NSapU69B70puA/Iwm+CHWG6x/DFSg
9BzXrScTdpuh6XLqndPLPAuGIQc+a0bQ9+qcEQdGsNAfrm8USAowzt3XFnC0YTwj
J6PEmdTiN7qStDT7wvWVjCTefUR7a74ZlxxDltBKyOxOAq55/hx/MsCEasN1Z6Ty
BzwSCCqXYXIRtCDq6lvlrGXJZ1Z3Xv6uJvWN/y/RW4tMJLABID43Winq6EqsWW6l
8707vGlhDgaQFOXVF4UNoIzNP2BJDBYWvfCyvcmqV2gz9k4j7LzCSCIxVcQBc36G
bPfAI/okP7CXrn1hL3FlmWBFugzEkofJ+9a1HpMtO0Tec0zYkW8Ck/gmMSj5wnvk
py2xSNMtmxiTWcKyrLUZZ7u5A5WFuc7LpHnt89tQjC4NBgZZqTNquPwYRzA3F0+1
wLt9bM4nVpsZ1/Kj5fxGAlXe6Tnv6DpMkY/8Ovu/oxEdlNNomsS35fz38I3MwcMg
w0iqIHqHYyNXDjYH4aN3JGNBDcE8yx3txQApBvtx1rmxCED9Vc63xP4EksjMIfyB
j0eUX2XeDAmJjkXwDJVke0bbBUFhk16TGAM7Fcn9PayiPey1SNiVKnX0z7M48KTe
rztBtlfIBZP+V8WVivClG85d294ghSKk+r015zokjgTOebdCPux7VFfEklcZ6zEj
BB70cEi37I8u8eLX/ZOMNXZWyxd72isqq4Cqt0xXAyjL7ZLT9skaIVrABpUKlLr1
NkDA/akc7SvDzUDprDDJuJiZMf+UxpdNLccRx+CC660YZccBQqUEnWuPMd1RkqFt
C8wNBr8sqIscwUs8c+952y4kShXg6fVpXoxBXZLAcZwomEy/KzWCLgzo9pZos2my
JciTMM6ij3eLOXZdM75yMMRCDKyDQE1mq/pUxYliHer3ScqafvT3eSojSX/4+wtN
tunvNwfERRPHhDHSsN+7Wnp8mUMGJyhR65yjp1op/5Dw2BaC/zBhmuwaV0feMr3k
5VSE2pVQ9K998HeYFZI2Dt0xK3JJ6nmLDbkZPzEAswKQNosbFO6qhs2Caz+FY84Z
ds9EUzXnpUy0evSJm7im3Bo61vmsU4tTqyiI0JrFDkVVlCSm2KN4jw0vHd9TZhMr
iLHs9VpI7WolPLg12qY/RacA+NCP9aMFDpgIMkV4J69sIAx2k2MP6lCLNTxJoAtx
LmLHaAykTakKrfISsgidVkc5/E6F3OuteNhsrqcl42Qm5KrxthaNozZ+spwwvN4x
WBeSU0Ucs3MamFarlfOZK6Teho7apv8kSkKBrm89MVfo8pEtzyTbTik1q/3k9ASC
paODzVLYNSqmjxJ14iPmxdUKrHzIywnnxond7IxpC+V5mDbUCFYSOULG78KekAEJ
0e4iGx9OYQOO3+JhCYoya6DpUTAFFtj68jXH57JY9Do1w5R8vezcPyPzIPuQPvxQ
xEUZVn9AhBp07O7JY8TC4EDBEGp3FI7mB40GvvWcKLLQhSFcvUntKHFc7JAb/QSJ
5t25hnn1tbd3vPtHQnIc1mofQh5nuupEpmS3GKFzpK7KyYb+YY59YCZ5UMd/xyhN
R0NZuk8JisCVejOOta3eSEksLQAarWfHklhECjoB6iuixJHwXZi/T4L88vlIPFfy
H6As8vmGG4TZenSU7ez0XyAZafB/z6TUDl9t0PonhpQNI/19Lc0Qr0aXZ5eNNhC2
NyAt16Mgdg+hHwRQ6G/vrLt9IfHF/LoH5xIv2Sea7fIOrHUJ2ookOPiJy6MdS4fx
mZTBMnAwHVGe0e+/92b6IdbD99T0B8DgJ8yitXfodd+C2oTJhsX4lRvfOwQp4S3W
hQEddlp2Y3bSl2xaTPaB2WpFKEZC7HnyXgjAoXvPede8D3ehVHqI4SuSGcIe5oVX
0DidnNge0rP/TnadfTxgDqcADwAcIqGFTkvpul/jMrp+4FXQjL5BENS1PUuiQCkg
3Mi+Q7qdKReNQFWUCEwvoY6N7Dyba+0mqv0dTFhMQcJrLhUu0FpghdDp1Sn4YW1c
EIYEhA7UOUCM9XqoF9BMj7YEYjitHvJc4ZpJfA28rBWVjlwzp+62rzCOHc/HUHTU
k9y3gFaNidsgVfYqu6kcDj0IBLQj2ZnGWMaEyeCV5dTMSl06xFjJfRmNpjLp4n8C
SVC0qtEzXQAeGHcgPI/zFLbyj0WtZm/EoEiR8kxl/prvRR2xvX+SR+hRmXJ1szLn
hxEv2Sv6opR4mfAQ/jgnRG1ooUM3FbUH2/tzwZhF+dnxr7sHIp6QuhOk0gw1TZQ2
TLcd+0dyZxFjxaocZIHE/ZRJ67QAuEuVbJZP76CzQaRYomK2w2FyNE0fPr+zsD8K
`pragma protect end_protected
