// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
`pragma protect begin_protected
`pragma protect author="Altera"
`pragma protect key_keyowner="VCS"
`pragma protect key_keyname="VCS001"
`pragma protect key_method="VCS003"
`pragma protect encoding=(enctype="uuencode",bytes=200         )
`pragma protect key_block
H*:G#( T'#])MFO2?#2BK\8_$1?3WZTN'61V?,11+9@U'6J:B"P;1JP  
H?Y4@(*U_]+XPG-*[9QC^:H=E4J05+:"7[+XJI@195- ?ND5LJHX?:@  
H*:F3NO&1FR7B2=L[Q!=+FP.)NFC]>N5%"0ZLS>DL1&KGJ9#OJ'5+"P  
H;R!\ZC<0R1H$-T+(9WS2+3^C548BJ.X*F)-_I&8"#^W,2T!'+B7-OP  
H*6407\51M HB\:J2PN[ .7?QZX^^V[YB<H+6DR ES4,9B19VKX!F4   
`pragma protect encoding=(enctype="uuencode",bytes=9376        )
`pragma protect data_method="aes128-cbc"
`pragma protect data_block
@.$YRS\>IBDD>H'/(837S>=0BW<YP^$G=6&5D9.Y9%.L 
@/P;/3#K<,<!<C;MV$G5JD,]/2J">]MSF 4;NQ'LUN,8 
@XTN)L*8V16_-1MN/D)EBM=BC$:##D:)QRDZ9Y+2P# \ 
@Z:9H_%U85OL2W9?#W<\GILSOO%.(<5)^&DC@H4:K/K$ 
@,ZO_,SQN[KKG#XN)9>#_T8NIP@#A^(8;W']Q]Y\.7$@ 
@%']:S=(J20KG)#U'<XI58>YW(.;@ DU<)C[H<<Y@VA8 
@W<6DPE<!),B/D9K>7'/$4B*NW"A*\GI5$>&FY0GSZ;( 
@"5AJOFKY80)0=BS*D.$=?R$E$&Y.3RJ:O ;$ 1_H# H 
@><UA3<Y*GE<J[Z$?C':.;.2#]2KY.241'>:3"K]HH<D 
@%=3OA4>KV^0!S<591)HZSUC%04S1^JG0E#S0GUL/0'X 
@L_%T'! W5<?G&-U67TI,M9&JL-A -X=^I>FLT 0S3#D 
@MA/1(L-@F*2B_0]#:RC7C%2G:A\$#0*./INB!LOTQ;( 
@!VB3?[*#MWQHG^,ZQP5%8F^Q-"A?X:&JA)P@GD%!=F4 
@RJ:9@F*8/ROF8+U@,="VU#Y@,10%6,KC\'*YOK$)4^P 
@N[<^&=37#,8"3Y/A9,-(4;\J9PS)<\8X?2+9^4D84W4 
@"9+,&N\4X[HW7)H7M+@SJ+[<0+_JB*;SBS8HAT+5<=P 
@2J=;;[%:+#65&+ W-&M//$=B!TTWB!IT_" 5*?=.@9@ 
@5FY!0J)/F<6&-MK&?I,EXBJ-F#YSO&ZN,.<#BE3HJ'8 
@YG\Q_OL6"0P=I"7TE$?J>,[ 8GEC/E&#7=+0O?D]MYL 
@1,6V@T&EKVYM_KU23*7)KIKWR;N4]C#>G!."%_BKO^P 
@<) *3<9ZMB36>E+BY]T7U",B9"<ULZ\=+?1RE7>&1MH 
@SF"VX^J"WUXU\YU3^_&+XX*__S<8NMU9!3-&5[N_;-$ 
@S?75R'#P_=8=%=]IMM"%5I$!?GS$Q"?2_7(_V*)6VEH 
@Z@D%\UU'%+80P/T2SB=BD"H#[\"*C>2'US:X6].&)YX 
@\XMC%%=9/)C)EA]][)M=P%7+\'2GU/L*7(],(.'Q%/$ 
@8_@^)U_!Q:#730>3JLC&GT/0CZ9EA)1K  [EP>_!H'@ 
@3QD(A9C3\Q!\O'S)&%0W$0G=I^8R=1-Z*TVD7+]8HGD 
@T_!B.8/#*6<U&YB:'9?^D#[]O;7VBXAEPDK:UZ\MKC( 
@WB;\S(4?LCDXI4%V_.IY7=CC6#MS")%OB7XA&]3OTZ  
@YTN@1J:PH8!Y%&"YU343R)3%G28R_CSKR2@KQ!CUD#@ 
@D"'U5U-C)/+Y55&E=1/.%6D81& -05GD%>YKDD1W/.L 
@%VI"HF/XH:Q;9?/Z:-RLB+.\9MDK3W..<7NLT^X%$J@ 
@.]%[)_5E'''2R%D5BL(@]&K$]18M*@!!ES<D4]PPY0D 
@LG\2=\(9$'\IJQWK"Y\002T63VJ;P56 <8J='A(P\RD 
@& +W#TA5H_Y)H 3N1#8[]AC*Q>4AXI%C4M<VQ(4DM[$ 
@6T J2'0?$JYAREWQ6>2)+PN<'(FB^"8-)'U;(AWL%J0 
@VI=2[V"Z+M6XF6LMD*UV8XA:^8:G!LI[@?ITX==C(N$ 
@\HU*H_3_PB.VG].PE;6A8N=OP2%YG\/6OW26>QTU?AP 
@GO=E^'S<O>+%D"*O!N9S&Y202[B/Z_G(YGZ.W8H":1  
@HP&N4<)TR38$WY0]9,TTRL^4%6%]2+?9X8?>*W9U1 0 
@0N/UP*S\VDDC-_LL=F6KG[0!_SR4+"&D11(JN7WMVRT 
@ </Y@.*0]?HCYU>1DQP^>\N\&NU;G/ZUK?B'0C=@VT( 
@QA!$HU7 <]MIM3NY#FFP20E.42.REP^>M(,"3<7. 3X 
@?@Y4$[DI*F&D??EC3A%-H@<U5[S8@)>'*^4#>V$Y\IL 
@Q3O'D$]O=$M?Z);L&KWV1-IM!9)0,4)-E%N-=C"1GW\ 
@,1!#)V:K.P[ L+QS94<3*3%>^+X<Z%]M5.RF#$#B49< 
@&W^57%8C@E:[A7B/.D]#LR'MR5?3T\<_Y%9&H>'4GW< 
@"W#5S:C?<=3W6=*P%"D(/ET%ROH8;#P(GC ?W$7)\T< 
@PU&09SHTS*%7F+F3CFD(%56#:A+8%NBB%"J"XU#0!RD 
@QN QP8T$0!E3GA(;?^1U%N9@&K+R-WP']+"4KX5_VM\ 
@63Z$PD.?!,X^F]*K1ZN:G7+FWX;&%-[28Y1&M#P[B-0 
@RW>X(&,]Y5B"71M!OREG^KICOCQ^()*%%G;8KL&E,7  
@ F2:.BUB1$._THZ]I@>(-98BV&FJ!D[8Q1TQB>VH(&D 
@_]Z(H"X7^^X!)BAU8F//!.4=D&P(]+H9J3!37H\(688 
@=6D"EPIX?L_Y[#A^W2'!,<0B9^$IC<2N)_:=E:BK]4D 
@2:;!T1-8=ELH3>'&<KATO0I3BC+U GK3TZKWNJ#6:S@ 
@\C+KIWM\*-7H8H,GLC_1VD@PJK?IFP)K>PH1WO AL+D 
@5ZCRX^DK:3JF?]\$6D++/J/%5E5Q8Y8B@ZJ'G<L@^$D 
@7VZI",O_X6IK,$O9=[=$-NKLY]E>S^;2S@O<;!7[6[@ 
@.<EF\=7L[JEF.H7-;1267H->9^SX%&&UERV$@O_E*7D 
@<#;>>D)7;@>J>[?I[HEKIRMEQ3*E/73<\UH3:'G; N  
@=/0!S:K>J N25>N+"&JBHK?M+.4#YC"&/T?0!#7R"3P 
@YJF5%0Z_)Z)NCASO8"?9XKB(CL9< Y!3,@8EDUZVB8P 
@][)A(Z;AV>V+OR>M2AK>N]U!:22*G\'3#*Z">\G$'TD 
@H?.M-3Y^=$5Y(L94^-_(E['2<<5@RTO(X$3L3%17D3L 
@#/?(1N0V45O9:E0&Q+KV-\FC/T/7^A<-L 2+6]9;1E< 
@.A\YK312##]-$D?*,O%=8WB-69(H=<LE&L>6U.]QC@( 
@6S4-=PUTB<;%?<QYGEW-&>[($U87+.4(+%;X?=;6N8$ 
@3O'XE[7C' L7EC"[IUCYAS*DDUYUWBX-!%ZDH'!%5]\ 
@0P;?17@T'^W'XT/!A6S_Y9G&A,L1V/WKYV*!%Y9"%Q4 
@&4QGM- R/TD7A3YG>3B)-$(4*6&*?"T):.,JDP8'[PL 
@LGD/NRK-X;!=8*Y*\^5"/2_-=9DR"8&Y%UJ.CAJ9,#H 
@=Q5]?*0'\KF(3.-#/C/+/X<)I+5MQ@F@KZYDB6:GWR  
@,/"4K_VY'#4$YXEVE*KNEDR[DDVA9K1("O%.("1;B-4 
@:#7F0OX%57BWB(@NI/JG)&:NU2_NACIN!%ZB\K(,.%H 
@.+PWQ9<"<N5I(DM4#,2?ZT,:S]#C6T)Z\4X%$LVH.UP 
@)/5/,6[YOL4V;.7$3S^>-V /$\$)6L,U?IVPA4MM(V( 
@3)L_N)9XL_D$X=M"]QL 5;ZN=UA$8?SWV.,/?3@E.%P 
@1.J?_,TI@O*09"&:[/\ZXVD0>M_2D[V35YD-!?+UJPD 
@TF$7,N@23(%.C"JHS5C_NL&60Q0!%7TJZ*.>@V#^(*D 
@4OUS6W%N?*FZ.#RMA+M%YO7W"3S+A79C -#P$IWBG+4 
@4QV9O3T [R^6(<>%%M&*EEW\%&EKK*,&PJ78)[<:84P 
@D'XKHU1$_DP9O=O1;'[3@:)ZK/7F]Y'=E^UJ17-X>U0 
@3I#U0:H%D0X+?;<L&6%'+?P/%*YD=T'Y._!YROZ<S=$ 
@*ECID;+U!^-;.JZW:X,\Y[@+[Z70+<Y"FM&5&LX[WS$ 
@H*B34 </VJ? &,//&\1D-B84OK]* T !K<MUUL[).WP 
@)H'&4&RZ>//7T],EN8OP% ,8YMW,W6028)I3O3%^$R@ 
@L^/8;5X*=AMYN>G@V@+=5@H"XNB> KE1312TYALEE'P 
@%DT;*(!ZC4)!MQR<KT2?3^. 3@'"VPF83:D+^^A5W)X 
@5N'($30B?!VEY-%#FDDX;QO&B, )D0* YRU[^1"[EUX 
@%F<ZYI2A.';.4(R;QQJ]4ZXT::MI9"8B/-;9NJ)IM@\ 
@ TFP\<2W%/9&FJ2)JRM\9,C1&JZZ)2;.ML]&5PM"7X4 
@(,8G+#:RV!L'^C)%I _7^?TW:/M7D^<A+S55G!VI,F< 
@=I9Q+3=,:-"TQ?,V@YZ:PVLKGG]01%^>*Q<#5Y&(SF\ 
@9?4CP]*H]$\I1Z7T]A4<\@W1MIX8CUK^*$]2D1<MF<H 
@)<YC=]M9^J /7^6(C$O"'R."PCUVJ)\/VM_+G;-0A9H 
@JOL$7TFGT=- ;G>0M9B<*+V%R39%53<1P"Q'$_1513X 
@'YHR9 <IEVR-2]-.IVJI@&Y+'Z\\!N"(\[#NYJLK#Y4 
@GL+SD 2#.4>)=I(;6UB=U!(AXE/_6GG^GBHF0GCP &8 
@H#0%R!#V]^,'#!0248M6-#94JI]V!(:.<MB<ZF)^=Y< 
@&P"W7N!GD/[)O\_H7@BGU3L?-C^&-(+(22['!/&"A^T 
@:F-Z9G,&1=]?6A4[,K8K$ H /AA3A2V3V8B-@TK'^$( 
@AB"@<GRR]-^_!SH4.BZJ2NWTQ#2_!L"EF"J)C/N4.FH 
@G^\OR0*\8A+":S6KP$1#=C3EH3C7J#ME+9&T'[?3?:8 
@,@(C=8:E50?UM4MA,3#KNO)B46IN1XXJ,L4;*??#A%4 
@S"W'?9&GR*%."]&BW<M3T^#0[PPLV04/HP?>7;S[H)< 
@>3O*L;,==9J)5AS%9X1/M]1[>Q'85^L$9]JU*8D6$VL 
@A*T'#SX:32UZ)5\I.[[^*;05<))D+DBR R$B2=%/QVX 
@<7YBE5J"UX583SB04)9YKB(OP_!% %#I&;-J_%LRLH( 
@JJP#_7K36#WA/\7L8;AK2D:@\$4PC!>]K*1Y/AW$06D 
@?\*HW)*!M/.+M(?3D'U3 ?M$MY(UEGJRH(U(IIG>W50 
@@G)VEO-J E)[ESMV9-@>FTC=9C%L[2.#:.*'X'=]P,< 
@A[N:7A+G&4BP]3;RP!I2VIB>\/%^]<#3M3B2GV9([]4 
@H:4XF2IJPLX[:CI#'&V*L]HEF,XLL( YI]^\QV5 ;EP 
@CA&_@X<ZPF->PZ9S8U5#)]59A1R9,5P$L*2C;P4%S0  
@IJG=0NWP]+6[4I$3@*ITVBD/@,/7&8#(#U_ET)/$'^T 
@R ;A@_&F=%9) .:9J[#]8^RRSYXA"8(0:R0WL.6+Q#D 
@+!"BG?'OGBNI9GUA+GN^R] [?4MV#+&Z4'P_B*FS.TD 
@^ '8 7]?%86O&X"/IR'$[AC'#.-9D .TSH2;&,@%X_L 
@^>]S]IN\!X/D;!I[2L?'$9QX]N<8"%AJF;[>V-?ZRYT 
@>7Y\W-M6074LYB8M&9N8)_N--/@_",(PCJ$ WW#1@KP 
@O4SJ!PJ+(0$3'=X2-4#FP^@\CQD#]_?X7,;A3$N$-W( 
@W,%K_@6)S<,5>[JO0KAK;CR_@G&1C@M<20.\(Q72A:H 
@ U8_K;$GL%+9Y;1+A0TQYJD"*J(_J>S?>'KXFAT&GCL 
@+TZUCGQ,51PZVKWG4"4:)P3['PG&.2'R<%C#F[%0+]( 
@5<T7=RZ)LH,S08)^M$G/DL]L2?_HS<1H=$V$;/(94]< 
@EUOCGI%+=R376CYY!OL["9&WP7%%UW2/ #%F2\NQ,@, 
@.^6)+:2^E\I\U)A05 MJ&L Y[H"Q:#1*80!(1=&@;VT 
@:XNZ]T!)HQ&VCIB"F)HHDV7ZY$5<PJ"9?$-5/R55B.H 
@4]]SZ4T%T-FH^SJPF1!\G0*C:&5;U;?I;"*=<\Q(S:( 
@K<M1."'"NMC?-I#A%$VL^"%MZ;Z9D36A,]#<8FO^H"P 
@1Y07R\Z<B>6%AY]M<1+@,'1I/<T&G3I<1?[,CG(_7)( 
@ ,B.EX.-.6&1%Y0E"MC&7:BCE;*(G)*DXEP]BZQ82)  
@(:U:T$\^'1"%]YFX6]!].>;?I#],.^>T+^]M2J6V \< 
@UL%^ZNO& QK;!9<ON$D#9.9FIA:K 0#8A_CY2[#DE:\ 
@OESS)Q0#!$SIBF%6!&'!94U-!*#=-A ERMQ2C)<>[)H 
@8'PVF;F8\U=3K<W!\,@SA@P[_Y#?6@?Y!,6#7X)&P\0 
@2_WANDM"-_3&1K=;&J%F(]/:1S=U&'E[JFQ"E%%S0%H 
@A]8DRL4V8R8-6OV4?CCDOV'_KC3(WLX(;KP5@-M4,2X 
@<J.3KHNBJ@9#A8U[#B7W%<^EG>@DF?1DD;&&;ZBD[MT 
@%[5+VC<4PA4GK;8"V=A'2O:Q'[_T4HHX%<^0R?"^^UP 
@6!8!]3A5A=,QS/2)X8*]PB9KH4OVO 5[EET*E6V-YF$ 
@;)Q:/8)O'$YV8+E7_/=#K*[)7X^*SD-_"/[O%5L_2!4 
@5P4D&?ZHB*LONRB>BS^7X-, ^]C(*VH;Q#,,5(@J#AL 
@31#=%X9586UW IG]1<YAJ F?YA@(8=@P]I,;]6+26-( 
@M/Y0P[@(UO']YP$JZH6%>O,S<]RAD2YV1FY&,W]A5?8 
@*XB3VY?"'!L&0URG1MM19: %%H(J6:K^EM$7$1$44]< 
@>%')MK5@DJ",D?""B<')9DIZ)-4_GSG;8_Q@5D4O5_L 
@#55#^!JG9EO-T+VG*#J)?*:W@D5/K-BB,%&99AKZU/  
@(=IN?,0+TA5\'IVG^$.1SK:7ZR!2#OZ+15/FG878QCP 
@ZW[6/3-V4H.I50+Y!03"#]OV2%1E&CVPDN(@*TJP0#D 
@/\X=$2:"7_^ !<)OZ]H_*2K@MO1S-CZ!+W.&%LJ!#"X 
@;!L3LEES1[)U#\PDP6(ZMSGODFXH7\^A& 27Y/*- G  
@$"-*$6)#'JE%MZU%7_"QL86^B&[P.!.M=5)Y2N0+D<$ 
@O7\W\H:#6PEMV!<PBJWYH]JV5?)2SJLYUB$W38PURC0 
@X[KQ?X0C!)L'ITL03K!U84%CP-Y&ATQ5T%W&",I:G.@ 
@YYZAQ8RT)@90DZO[='>#_TR"L"VM;@%L>SYN2TLP,N( 
@:Z5G:P5PKV9_[Z2JH"C^/A3-W"=]DPS1YCZ!>$LSI+4 
@"<"BY0IG]!<FUZ, F8$NZ8RZ@*N48:9EC\&9V-Z8Q0\ 
@_3L=^)5,DS1HK_\Y@W@P]BTPR#I:&^@#@]_;32GR6KL 
@Z<4!+#A^0]Y[AWJ?_!+@04.2DD)(5U9C(.\1\I8RY4L 
@PTID5\6,=_>!]BQ"V1M*U'%I'N#VK(!OGZ/&2A>A\G8 
@>G=V'C:RJ2^.L-IKB3UZYX0 =Y[O]4XB=^F=DK_(P>T 
@U$JT7QZN%=C4L"0Y7FRKA0W6BX"PR7X70<"I.HF0-&\ 
@<G.P\5&5Z5&RF%$DD^==K%-(M'Q)Q<VWM!\WQ,P[OOH 
@[PQ&5T/+5ZEF[ $H,C8X7>5![:19Y/HJOJ>!%T_PE"  
@@'TB[="O&U^8.))LK;26[)@L$Q#$) 4)#U0=U%( 2C8 
@M2?H#,\=6U)RIK[X%86$X$ZV,]['RU]OTHFOWMRU20\ 
@R00!77P?E87<UWN+,4OX[E$(%W*0%:=H@XJ_H^E,R#< 
@GAOZ!DS',9'M)TUQP@I!!/!3(>>S!-,SY^=JXBFMI$< 
@&.+Y >*QMU4[//B(\7'#A]O=6N#]06FY:IMZ7',1,N< 
@NZ<WB7.<48RU"5M\9ENI9]N?H;?I"[C9"&4$*,6_'H  
@"),L5Y&R'2\"V!NBZ3_P^ST_$\_C(3F_D"K;E'^TCOD 
@*[KN$<^]B/!$_%Z'"!3Z<,<1@6R21*#\G(JMR=$?=!$ 
@(+PG5:EQ^2_-I<<F )C@,,YLHSD48/**&#'&N91"%5@ 
@YN8?H/*0=N%^>6<!HA5<+IRC2L%5,X<W"7\?Z3_]$^@ 
@G^<!+NORWXE]_L?[XXF[\_X-@9I_>NZ4)?3^J4RL*SP 
@?N94LLPZVNTE  ,MR'U5G<FS=]M?<#)T#5A-;N\.Z!P 
@56.<(ZC:ML%D<H^^]]J^]1>G/3SXO)2\0%\<8#]6^UH 
@J.*N9+MZ/RD*GJSU*S8M'!0.%D4DLBY\O'"L?I)[D5( 
@54?F5DZ7Q-&RRXS]>R]/PRD6W)/BER8C3Q;(:1B^O_T 
@Q<.^\_9![Y)%?S$JR4!2'7XI[S)N2H*_(N$V_#@X=PP 
@6HH>H$U( ."C2G= 26V>@F?CSNU*-K4;/GWU-\TH5N0 
@8=GA+6\&VXRA@59$XR-$D&T+FH.C/W\):,E,1ZNM<+< 
@DMR<4C*UL)[7!8$!W]B ,X) >VX)2)TSV559T;R%](< 
@#LO"*/L-RX0\Y6'LXS&U< V_%):S>H^(:!9>@.S,BK@ 
@^:R>8SK,G)ZU2IK^-NR)./8VG0=*H"-PV6/C]&^WU.@ 
@(BQ!=?VVC$.Q_^B/5VWGP12=$9FM@*[F);9%,AQ!;YX 
@0/)C5>VRR<4A6\78BQS(YGOG6 %UKB4I_PC^>YVS^>T 
@>\_NSO+;08P@=;%H^CUI R,G>"/'O"I%^%]:V=;X4<D 
@.'%J2$",>&HV9NU0IET_9<#P"=B"JPU EP;R6BN8(\0 
@3Z"L8A?F -A 0C=329?H-&]O'5\XP?.3TJJCW'<-)A0 
@/55C?19=HYW[9AX7/C9YR,+5F<*$1RUZTB-#,*_%]?D 
@?1(^&><G::HG(@P6@V?!*K4+;I_RZ)OBW,+06&\IU"4 
@DAFI<$?I4:9_[!LWAL+;:)!EL0LM<3WVC"<EC+=2=ET 
@^"/[+]/7L]IA-RCE,<EQ'NP8#3DEE'I)C65;=->4>]D 
@8$&B=$8J@.Q*'6;0_J$Y5+6F0*8HYR437M/BPM@**]< 
@*(<9=IW$( +OCGO0CQ,_LG!_]&39>Z)8*"*&]D+@&L< 
@]6[E\K=X7$U)MRS @IY8\D:);;JTR$(.I.'WB"W3840 
@B4/##P@Q:C'$++[LDBY>;?4_R.)T:"]YNH^:G"R=@,D 
@V2)30U)2_0SMXH;H[8)6-"6A'*,@+OP0JRYJAN\<5"@ 
@('U6_6N!/DU.?*6<B6TD2MQ3,V+5A@9:$+5\RL9?(T0 
@;CK<S#BR&F!D;RN#[R@A(X[-6N549<?\;YTU"G&S!L\ 
@T6%9[97Q0&0VNH5U3AO=^ S>]>(@^RXMLKD\,7,@C;L 
@5*Q[S1(O0Q7!$3;]E[\LS+BY#;FXH7V8T4I1&I@:BFP 
@VEZQ+8&O/"-%U)?N FQ9D$BX=$25&ZITSK&";5P]+3H 
@'3O[:5NQ!.==  6<WC"[H=2'IW,P#5 $;X0"0B?R.-4 
@1ZWD36Q.<=V9%M^-Y[;9-N>[W%G/H7-K8:!BNSZ5Z9L 
@2D]:MI1/_7F^'OWQ^WVR% NWLWWU_&LK*6;-X"Q?,7( 
@:K/66 J*U) 'JD516F$DD>+*JVB&PZ$Z3X,*C*(S\8, 
@]?0S5,II[F.IM.4'2^UXS8#T.OR<R]E2%R/@J+M%)>$ 
@5BVR9,#BU41>(Q,*Y.E-0SUV4\#>/>K%..U0AJJYOL, 
@J1$!QG %.:W?1@690: J+.S"#*&MR1L<Y%+H) 8H#)< 
@A5WM+"!LYWQY!9):+O<>&=1#;WRF**3C@-IL78?S /@ 
@,6CS+V([<RJUVS,Q(P1&%Z->>MY+\D3,?$ V#_X9E(@ 
@.E]=C%B5D<&^;NIR 3G!Z\]1-^+93AM=;2)SZ"6J*AL 
@6##6+-B@M0VVCJ3O"+IH[RB*/G+O#=Y>Y[+0_6!Y5$H 
@\LBK1OZZ#U_15Z_;R#Q+]_8'[]W$][\Q7_Z^ ?QX!E< 
@J"F<OA%7Q;,\!S]]P&J*UC4*>E9F&>?[/Z"-<*00,U  
@G,PDU/3EE11MS-.0M"S.- CI?X!8 (XX._2\8,(RKU$ 
@>Y+B$Z!4V&ZQ3#*H5AV)+73:D43W%8UPC 2^H;OZF>\ 
@T$6%2 )Y@=W,RO:]*S,MO ^1-,E+R*KWPT.QCN>BW1T 
@@870K=V.JEB!F%IN&?WBA6%G_$\)UE+^G4XT?UH=.]H 
@)=9+";VJR3K)BCI.M^CQ[W] "GK%2^@]?)>( AUV,(8 
@\(IQ=J<()=^P;+PPS=:WC76F%GW8HZC%9C) %J]U(W< 
@Y)LP[!-P0DV\H6<W,;K'4.@CYK/14R<Z/G*LC78^A,L 
@,>>$4X97  X,,U_SA>7+/2;A#(N>,#TXQ"@;GI?T'!@ 
@-LIC>]<%RF<XXU/*XF]D=;)3QL6F-]9(^<76YP:DU7  
@R" NW:4\AOT)+7\.ZKQ=OO)^W_K>BHPE=F).VKI1-@< 
@FF(KT9X@C:_-XP1*>6F'STW-C*TW3Y]UZ-4KO5D!OBX 
@S.Y"DKQHY9S2<F]3G2/#K&VC_7@4Z/6L#+3&(C<HRRH 
@]5SBV%#Y"XI.S()J+& WA".*U,* S5W=K"D$@%K5*7@ 
@^/S\M#UBM+L$-HF'3PB4J_5MP!R":2GL<+\A%;;F)X, 
@DP]S5:(1NUD6R]W'L?"G4Y M1]H+$Y\B4)ZPZ3<@HPH 
@)RZRT2"'K_S#/3,@$BF]V1!(^ 0CJ39NH*C.0W$'-$\ 
@L@08&P?/%\\&0;S83X:).8P]F)4M<2JKLC 3:OOIZHP 
@Z(@FN2R$Z)Y4.-=NEKL?'FH^):VU?.\4;"+1)OJLYTX 
@!3_! ;,V++T6M_O-R_6&D;T]W"ZKTK.#&L6?1$R['P( 
@*4GJ(("+X D%M1R ]-'@RA0]HJK8HI9YNNV.4R_KR1L 
@,^%:,L#O5++$<> "UW[F-5Z_3G>),I>#&VR,?,;&>_4 
@%* 5.I"0$)AEYNNO@LL"P[$P.;OW_HA0UJTX(6 4\9P 
@U5"Z52/2AO1#X(2C66C,OYS? .2MXC66BMERD8Z4KA( 
@6;:H5^&NQE7^28(<2K5]=\NSC*]W(%\:$MQ]44A9^AH 
@HTIJON$H6Y'Q!G2!>+\P)9TJJ8+AW7I\-/+=#C-WW80 
@K:7'):BN"GJW%DJ,A H235;?=6,(@,H!(+DA+I/KR<P 
@=CS?_8]-$[+FG6)+538C##4((C]J?)W>'0WMBKD1QMH 
@G?TBKZN<J1L0FJ Y1PG%*F*N'V(M]5L1FCC^M/-J]J  
@JH[F^:7ZZK;<RN7 PZYE?2*H2!<O%]T"3$41WPT$Q_H 
@G)W+VS?6<AGZC1T2&@'&2V\<<HES-G<J-9H3V.212+L 
@JMPL:)H%I#FNX?M\E3<T/9SN81 #=*D8@K9:ZSYO8S( 
@[T=>%V^B\GVF]!G'+FTW4\XD1E._Y1=\/<]'FTZ@,HP 
@#X*= W<0/%[U*@W2]IAER/>E![]>R1Y(0JS)O?O?OLT 
@:!=:+B-G4<S%DF1\U7ZE')?;J[W-X"H761(SCJT580, 
@3:ZRU[P)KX:2&"&1J%BW#JY ,Y/^U6&=D739M1A8LHL 
@KPX@ZV9[/:2P7[S.KEW$H"NQD[O4!1S.ZZG:X1X28,L 
@TK\PB1-TNVR<-C<!]Y<<0KW^N!D#^VZ"JL9T=EHJ3)L 
@9HPY#GOMC(LKM_R.H"(@B\9Q)+[%)UE1AB0G[TCPLGT 
@=,4 S-FSQCA.ZC>8@BQ/YW'V?TH.J+-Z\)[I5:H)%5< 
@*2LLV-6BI89L+;6X<>*JQUJ?[L/X'["&H.T+%$II./8 
@-EVQNK?QX+&JQHVS"78")28\I,&"#Y3]LH&B-!&U4:, 
@Q9T\T"M8(WS%>NYHH=91'G@-QT^-='  ]YZ]4#7MJO@ 
@I ]P_8X>_>+E&7#Q)_] C7U_WPWBK<QBBS. 4O-A-7T 
@=5T'-J@VBU \?Z[EF%G*#V;M![F2HN1^^0(,;">,HMD 
@2#J];)GQ()I7?X@B^">/6W@/D;J'AOI_TZ)?'6'IR=H 
@KN8CQD+^64 *$<,?EZPJ']?^E3K9RV-D:.*34F;T*C( 
@(#)L+=E'\F^ #N$SOS4,3N?)L3N;^*Z &/CN[7:T/-X 
@*>)'R/@>/S>%"[XOSY4/^\,1*W)_A]28^BVF]@J&UI$ 
@0R)P?]T^#T)W-&* ^Y3$\:K,B5@.?F/; ]HNJ[GU0+\ 
@%CSI-7L]'JCJ%GKAEWJ9,X^">XRN>+N'S ?^<S\'2:0 
@F(R>.,Q*4><_&1HC5N;KFNN4H&#CA-K==,)W;H#0(ZD 
@%=4WLX0,^!EE3 H >QLJ9<"D^OL#.)TDI^')L/[QUZ( 
@$F*1QGNZ]>'DO05X6'$?+(N+!'3%,+!=2R4TF>(4BJ$ 
@M$[VAHPHM80(>>(9Q:CQ#2_KX.ZGFAU3_FFT=*)Q?O$ 
@$^F33+NFX#4!7^WBK4Z.BOV*[@,<\E:RD>&2N5#ABOL 
@8 -_/HSUNMO=5Y978'!"M%.^/2*%:?_Z$2:W+0K*ISP 
@,^LA+/LPB;*EH!@9D1GTZ4D*3OP&X(6SP.A&=8R0]R4 
@=D(E4Y<&>JI<E;JU%IVUL,C7A\CU-Q^0=*$F.]5G4M< 
@?"P$5G%Q?7TM^-9-8+36;.IZMT6[^QXWO2%C>TTK_W< 
@SN7%N^D)[TB@?1RY)+_1A>5V);Q%6/SN]++ ==;D&)X 
@TB-O \U<E6VH'^_^M#2!"RB^<',#OETR=7W(45?D:U  
@4AP)K2 >@QF\W!V<DT,:=[)0F=#I'/=2P&M%5NOB^+L 
@ IFFV T9[$QY47'D&BWHS0J?*."U,EY[B]K%7T9VS_D 
@@+EUAKO<6=!71Y]UX\>.WX&61.3I]R\^"1M:I;M_]\0 
@8.19H3 WZFD;_ZBQ$T!3VEX+>?X\7M#_/R:T*J'HR10 
@C'+/,K.Y'G\'$"D7-8 8+/@G\ZB^Y>VK):)2RE(?SK@ 
@F"94^4@8?GYT@.#C0-13\H[#?,F8*T8ZA5^$ZWBN8!$ 
@QUJ_ERK*S$".D-J9)-X^^N. 71L]NR;XTZ<VS#UH'3, 
@B%R4Y6:-?!]U%*-'E+[9^A %,;LO-A<IF9UC& L3HZD 
@$ G=UR#0]U*I',(]6R6 Y99=;*\T'FW2Y#B5EWQC&8@ 
@[R7XI8A/(7.:,Y7Q%PTV8<549'L6'EJH%T[T^M-WJO  
@W0:"OZO,4% )"\F!4 %WTB#1L)FPSK8$9NJ0!Z"@M<X 
@%[6SX!*PI01SE5L-&#V+QJ6[FHZZ_7$E/)24"?%/F*T 
0DW!S54Y)L/^1;<55P"]K,P  
0\#/C(-=X84Y?,B?B]XXM[P  
`pragma protect end_protected
