// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:54 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
HAAvnHEG64mOUcRHME8RlWZkTfNaE/DnKXO8abgQ/0Dx3f4Xlugdur1svWJFYanm
OnWefeOeRPZ15HsAOPU9hzlao4WO9ArLVEmVl1mfkQZsJ5MC0DZJEyWBQ7Z0N7NM
CW/hPwMoqWRhUHT8ghWfWwooIPsgFkZTZ1L6r5PJEIE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8016)
4A+Dss2tnZktwqRFobqVKwwH6Y3T3iz2vevff+HEwkD3fZwlb00b0HblLPgKwxne
8D0KCrSDtF0OfzE/p7fJtbbhoyPqayUrmTXmWKT6XHWaFbEvz1aaye5nu4dX1vON
wDTOUHckN86ePe3eHQw1rIKgWKgPJKXoflmVmyRn2e2HKb1e/pJD+8A0xOQ9KKOa
C4i2gNSmNeZSnSq9YoXsmw8Nwj9dyKkvTdAJptGQZxATuwebnT+d5VArk/DhuhQW
IYT0BOU04dIffBeNYcYV15/VpsKCjWnI+gpPCWMhz0m9keI4yJYGDWxAYRxD4fmx
1hYj+OHaiPTLTgpM19TZ3L+3g7aqzcUIMl1kO5+3zghuShvfjHpcFvkSya0mCnSH
lTuiMzDWvMkY4RAHvBagySQfo8l4mzvU1oxc7kdXYhXicsCwMv5BiDrHlSVAFl7k
+Bc9ELqLVHNjq8c46B6/Kk1Z8QVK2LPRdwEme9kOWSqtkweshOWqr2BuBrmd6Owd
2tJTSvqN2dP+onjTGYpUPzTBk++X2bvbrsOVaqxi0t2RGP0NKe/Wj0K5UZ8gNeE2
7m0HsKv94wYiPe/TZHFT4eRscSmcFAufxQ2dRYBq0wxviTTo4TCOgj/yXAvFIfXA
CU0GrEpGphD7ikdTdLL8s5GFPZT9PpX5vkcmlgqn2enlurKgvOU2QHwwfzrevaXZ
wPbYWZ6ypB9DyBuzPWKkQdSh17QY0XG3lwovD6T5jdYWUyFWX6XpaATF6vx0wVn7
qqBrwebwzViEQ8YIa4sZT4pLN70AsNmaRcTmnJM8sfWDEujD3SDUpkz6/MNwMRdq
OO/UVgD+oY0KUAvDoWHG17egCsQhP0y3A5D16ZnueZWNcXz9pSWuQjJLoZtx9Kf6
PPJJP54qZjdeqoRoVM8P6SGcCcwDYLFSz1qlhIomRjfDwoXsJ/1CaL5usclzQ8pE
hOGMI9teanu7kPpJERaxmf+ssnWc/3F5KU1/3LaeYz53NV+yTYtiIILfisP/Zk/l
mEMzJxHQnZXnPbDZpNEljCKYUiPZubHbQurOZZinsaKQIcL/1UyFfhb1c64ajoss
T/UnPDpGyFRIz0z7mtXxChnwVg1+mQF6NGHcg0SE0nauNruO5NQ1Dhp3twdm9q5F
bD7ftfhjCEGEAwQK6mfvH1IoYx8WjxVmo0VjxeAuDgGojTNz+8oR7DxgV7u8Xm3E
PhfuNYuNWKCYtIVESIO+RtyV+5meZAHzNChbNcdW71uqmlXY2m86DzNUOJ9xWwVG
dtA8ZJ5XBB6ioPAwQ3k3bPoU/CnrsdHw7JF0nEYdgvzP7RcsCqQwVqWpeFL9GP+2
j0rlkZ07kzefATkmn+0ndFsODc8ezWtl0SOmthZ1NOQaNrc1YcmLFNjQOph7mSLQ
NIIUgwiAN4g8tseEk3ceLiROtdRD6ntpOT8rBU5Tj9y9gGpXRqEd/cVnvNs5idzb
a71Noc+c9GUOJeZy/k8x0H/TCiwSO4P/CxVFhMEW1D0igC3VaYwOUAmacrC11mxY
RwfvHYSkJFCJwJrZPc/Emc+JXfAo0YAUh+YaJ51V7wRcIqW0VL5hZHd0PYBMnVpy
bZnPpfe95vS7Uhd3y1VjTPA6uHn2ORm37ZncDZpN7F2UfDFttY7sjp7KEhfSV1gV
eIkAJhu+b35fmeCLfzGL4aQjVJGWVqk1qGeUpKI2H3HpSi7yKcfVGygyCHSvmJSM
uHsO1r3NB6BqwwEqH5rd6dY2MQxF7xGNraFzYUeS2E86BLfjLISQoZLMsK6msT8u
wvMv2rWJ2LM3M5Cg+gKfbkM+wnbIptenCwMiX70CIEtqm8iEZBgMbXTuny2v04yh
Uz4IfYtY8oWZ0K2BWvTGjPwth2jMxa6vLu1ecAR87VfyBqD2BeNY3e8Z3fPOUhpc
6qxWWgg1Xzu6Yaw+mVDlJ1O4+G3HKKLNnV88vgWazl8ppIVjsX2/4BqMIxlIBR8O
qKW601t7K5NkzBgYGjhSriO8OXEV9qJKGojIr8N0E+DoXId+4AKeRMkED/6dog5x
OHyrtBVeq3hCyxs6Zk211srPZcVNYW1+GBFg07MHbyOU9iJm6TVNui39tO4uDhJH
6DLbhDw4wanbkPfRxhc1YiLo5jwa3FJOC9iNJJ1Z6je2E4xTn6pqkALUpF8H+f7h
CNHjjyqwzIaDLukcIEbYJTLMnI+wv2PZRfPmi4MXN/ixAppG4EfF0aeT2CLPiaTw
WpX7IbJHxu/0qEmazvI0IIcjfgFDLui2F3e/ptcHTLaRnf5yOTy8VpFYEQfzNUIO
VDO01rex6Cy9417dpEMn1mBoBFoQ63li7XEZWdozgkFJVj7SxEqt4ZrIRmAWBIiy
Vn4ok/sBw3CXVWuQbe8YB5rYz6q5iMdOSVeLm/1cl6cF7xhJg3YMa7eKiEwLaZth
T+U8Yslpb4YZ9YqeO0bk7ldzPwqBeCKjFFCx6NVcHFPgjEkAcLT7SNzUgYr+nwVw
ZiM3zh+RpTSSRNUNWo4kVF2A2UXTurNU5M2AQ9B8hoWV773w2sXF79VHd3r29R91
vY5EWZEwqs1ZJLYsG4mBFwxpX82D8ETX1CO5hQqf2v4UfYqBXDe9bYYHQ/4UxDU5
QkMg8T27gGAIa5O1j0cbTEvl1TTTkdygJK9bNeeQkeLVUa8G027m/CIO91p3WAsh
cizZy5WlxBk8cgEbveTrSEb5FKrg7yVbjgeD+KLuqh86P0HalD1NZyO0V0JKqlYG
BKku+nNmMbHKZ8pv2uAcLEw6xKEbNX97WwEbNYZyF3YTlDmEqALgFUFYRDF13MWN
CsHzIyzGkbxJv04x8oU1RSnpc0LI6AA1JkKoK8BBMnNmacn+H2vcTV58x4HV99ON
vwCbVMnGw80atJHPIi1IV5QP++8O71dgaYPqqjKZ8GnQOxIwfMlXT/cAewiVUZ7o
+NkgWf4rId1J5SLfEtwBjVBkRQcg3jQPThEbN1wM2pvXPUjx0V0z+OpnrDDamZI9
8gHvmqmfgHcGG2+NzQrQFpBSHK/wqthbkQMZWxI54JTR+D9WbmIPlxQpbCR3EjoE
xfnyc0lmDwA3mrlRGRcuQ8V34KKt6cFMXuKwewmMzss/QNTC5JHeMmVNexSnhdIg
bvod+pPHZt/6b5KxjHrcvg+IpeMerR09trp8e35wYuT4YL1+KJHQidynhyQWvlFu
CnQMuXsrMQNR9b7dQ6GX/p8/gCfUbGx1befi5z1SgGgGG1osxcEJcX+Sd9JL0ZjH
fbeGF+qS9stN82KHhwav5ejcB+hR9/CdGD9+gxGw4I74V9tVljMqqxoa5MR9PVDQ
zAtckeafwWDVfK49urQgEr9Y72KEEM9YAzQoGc5SEj7Bcu/JCxYPdBCjkL2DikU7
f/kUnpG4F+LPcRb4LS8zvwgfOOQoAiS+VLiETGImXB91wAE6UbUV/bZ2sC+k3tmW
E9j1UMCMzpaPX4yp0coLiL0IiHQz2a0JQtKKAmVwJnQ7rgTiN3rLcD2YmCGC+x2G
ZfIsdoyUlK2MDLwvW37dj1k87m+SpIffAIzBzlxfkA+hQo1V18JXMKccZf344OxZ
UhBjJSO0GyTFOppD1xf8UVcOjTzNEMB0s0tiOv0vdwdrI63PnwPDSu6GgsYic1yZ
BZcshaeDLkrUsAdrLrD2h8Koi1YxiCUPUqSXrUAdZ9jFS7BtvcMEHNs3ueRR2ydd
5xx9l4CpURxgduiVMgYzE6yT5wFnfQ/IGHiODdJMWOgJ7j/pcDbXiXDxrGbEJjg/
GaPz4F0Kc3Fp7zP7sMySQE6Ym9CMmVkCI20uqSQaInhlKKJaQG3DLJ9HZU7/M5GI
cDxM/MzXFCEcOkLEl1iqBlMYHP0k4cOSFW0E15NDrzfseYq+BQgLhGUNe/+z8D5/
aAhOv3T+0umopgHpDqsz00Ao1q+sHnzs7BsWzgKjw0Xxi172iSBaX3GmGnNj8lag
NRREKU+Wk5Olq8RjWoCK8IGxmxYk1CwONW+00YpydGjS+bvHtmB5O8HYZ3ZR7Iwi
d3OCssg7/CljVjied8Pu7NUfLd42TM5sFPkw3hnvmEer61X1NJ6g9N/P5+AitzXA
nIayt6y7lZZqwY4k7fe8ZWGSI3FsSv03rSPT62EdeZ++usmIxq4/ldxpZWT2wZJH
tFvOP3iXsIgm8JEiOjl+Qn8jirLEXYiHQBG+8G2jd1y6X0DPwfv5bsy6m+snuHmQ
yVyO5Eq3sVIo7qal081daEh6jf33IN48Th3y6U898oPNi4uPa6p9FfB0ia+WzmDf
Hq4EX9OjNBnphq9HHWwXPDmo2aXz1NMtq2eIcomUmwf0uQR+GpTZ6B7qFOhEI3wo
cpgAIx2HsijxtrG2oNHxjnXznGRdYaj/S2Ux/wX08YanjyvCJxOkZNT6kEhaj2x3
7PwJvuX/xVXNu5fVso6h7EwWPNGHtbhdxobdDgZ2h7BozZKWaeD1aGciMQosZ0Is
G2wvW7/GnmXouno4AOHtN5tns/IC964gH+8xpDDZsSbAuncUUWsXbqjc8eiRRS3B
uB7wvWNB1ozprqxvVBe/z8YyRuPd8+E+zJmjGX9anLZ8SjA6LrwqdJol/itUxFA2
JA03QiQjx4Zq7nJV/yIEYHYFuQb8DzQZbtqTzN6iSTAqn5fdckzuJg41UhIRtXZ1
XDz14ieI1Aitp23iGQx/qneLJCDcc7nWwm63baePopSTnsqJWOhn5O86XADzTzca
ifoEKnlPISY2no51CnsJxsPCGV87qX/Y56ObT6MdtRGRIG6f1IyiQ615Pd5VMtUM
6eyfWmShw24nxmcP3nPt9rjs1F45ZOh1nhfwlL3jr3e1of85aNXRBVX4CQAYmZVZ
1CnMBQ2bd5wGn+zypHtGyQ3KGJ8eBqfwxOZB2lLSMS4o1G8jptv5VxACvBSfn7Gb
IHbdOB1fcrFyWKiMcC3dPPT1x0aRLAMAu5VKQBeWhj3V7YUWFRQthL7li0aBmzRK
mhpdMwU/LknzCsaNZKllhST6N32UB18kq7zzFP39Ia7w+e6UXdf45R1lNBqrEaX8
1OIEnXjCAZ7YpPuteMwve9J23mpKNnLs5QnOxj3WFHd1Yo709K9pv3BFCkuy4WVg
X9SmJb875WdPiVefZrBou8v3mAJISKO0zAMfLU3GTKCi6qaxFOHlE8rAlIFWZlb6
dqyaiesRYtf6v8uxp05uDPqLQqnt0jKhQ64/MhVMcl1s3edYFiPgC4Vosx8BwEky
wqOfA9wV3Jf87uRvEgCZHDIIfcCmZ1aIBr2lHx0m04sPBDK7axV9NIIii3AOcSGD
Z6G9BaoTScZJgwhpF1JR8xvKEqK6bTBkFPX5LIOPQShr/R4vvW/0jX0LFi+PTxYT
HIWOLOan587loKGfcQDedqdBdcbJj879uHssrft/Uk+pkwbYapV5AAbMhPrxw5lV
Hb5DDYA8ZhEj/w450mkDi9rsoGJytGXjPaDxZxULfWhyBm+Uwzcdnqi0Znhk8Ht7
Y+nvIX26ys8MUWLUIYI9Jt3xKkW4MJZTtq14G/aZlLoPi1Drdl9jZSQ+Jrb25Qcf
AXwCVhkisxmHByp9H1YsPZpCskiRZqi+5CszF5JvybteHNCTyKQZrYk+8bZaGwsx
H46SGJiEdVjfU8yelU6mIO+5JLqGmFFHaGvmmCnnvJmKMgQXPcrbBjlL8i9rX8Fb
Pxfe/T/F6tfzdOJAwLdFb69wjU3EycvPnNlnP763N15EnG1749oT+lJxHYXxO+1V
lQ0ScYAOyEP9NP5HJyLrDQNxmtx5DsNJXKiNuvodQeIdqBGeh+L76nbtl2I6sEtv
w/lZj43VlVXAk9lwQmCpBFeTWPckVe7YqD+5h72xFvC7WA82QXjFbyhjji+dxmCL
2GVI+yESnu3X52r+977sAIUtQUo5/bfesxVheZ4Rr9O83OjWp5vDtcyBBwSVSgIE
p8iWA0nq/0hZ8Aaj6Fe4wgbS2Uma6N/frIPcfGuf1Dryp+eXT+xppp0GhW7/dMww
NoHZhiWO02jELL4fjddMAKyYvpxEhxW5F7QUkrzChIcipoPOqm8guobxAT+6BRS7
TDAaoQhWFm4I2yXSCyGO5jq4XdBP8d91LKxbsY3PpojaZXUSwkzwuo6s6pV7gTG6
1HFyLwNFCjWROlvQ1K+m9CjOG14PLVTjSzGxkE1iQz80f1Wdq0wpFrED4XsBxAyf
OS7XAGgQQYgy0aNSEnlsFRmpYOw/u5y22/S0lpn1oJbiwNykUKw3uQJJuzQ6XE1b
Cl6f86cDusyxTV5arKeR37ujO86fpUTggxfZg30wWMzfkdE5VRQR7S8eqiWz7zeU
zxj7aHAnNhF8Hf7hDmrK/fh4IAxrLOKdxUFhwjvRLw1rxxxg73bhcZKzwUWi6ahn
7k1RjMMQT32WLndXozzFnh2zdqpYtlVk0q8wKgt19OPmcwjeULgCHwelWfmdxfhJ
GCakpp02boo3ZJyLiRa3kYxC0LnGzoxBdECabMRR55lyvm2fcFse6ACpZUrOXqwi
RCb0xkZ4jETA8Re+1gjz+GYrV/b9RTYRqHJKCafdRq2vUachiVeHQC/14HkwgDsN
nKLCDkURHwH4VQPwO078RW29Xmt0G+Qjlw+sOMDOri9pCW6o70nwuqO3bAPeyHoX
Dk9LrmaizloNVcKRMzwvFPlV/U9w7PnjB+/sqL3myMd8ezizdfJ1GzWy00tTfrt2
QipIuVxS1qNbXYh4yfRqrl9va6Xo2Eg+v38ePVDTkS2mMfyn50lAQ7hC8U0Ub4jU
Reja0wDwHgW8btJSrolIMMH0T9S1yLwCTGo+dcgmxMea/C6F20e4iZ0IWLFsXjU3
TOC0IWZn8VBGm4D+exqaHYxtGSJwQMLFOfV/l+nExkjGbo2eT1wifQs8gDo1wIGs
1P/O+kGIkafCX81wpqmzgRdKy2cngpCeHkMeHL8UJzLD7gTiBYINkMn09UnsizPN
D+HzBsImS1uqwkzUZkn+l+vjC4LWB/5WIJ+MwCJ5trwgM+inKNv+wTRJskmu0sNj
oXpO6QSJ1tin3mFB1SES6Nn7cVjBktotjxef96F6PGY/3Uxp5oOyUSYuNWQ+HwHs
7ITuCIYXrf/Y6XN+6E6h6mvGmkkj57pkuBo99bRZteuRd8xP20/FzIIinACg+JLb
L8qGYn+UNnN8aquu0uoRBohWuTr15DvT3/+giBXzmIFUm732qSkQxYQzzIZJtueL
MeJMnn3gPLUPo+xB7GuCVD9D4hHEfo2fC8XpAUzFQJnW8B3CaLv22wY/wHM/oxhJ
G259BlwZHPhgXOcL6B4J6PvLoYXCewAois5/updBn15ayxzcTxGSbygFQc8sN7lm
gPAOwa0B4sXz7AI08SwT9Tt72xynEHGkhQXN53+MEVdgfhGaFFw3kUkgeG8P1dcQ
mr9hnItORbjIxadu2t/tJm4ZqPwLwvTYNBt9KYOoteVjqf3v+w0HF0PqkqB3i9jI
8vYOQg301/DF3NQVPBrqXghSAoJLzUObl57axx+wsVzqHsKNktYvv0MWBq684m0T
aosoOVVaBax5mWaYTJRpYYOCWVv7OPTOanxJs2hAcD1SDbf5yB+iYaIQng614YzZ
qUFyh1DOqfbyfDVx04LeHcHRgdjLjpuuE65Tw7N3qjDN4GwwdzADyKMvsX7gHDJS
Kn/b2OnCYMensxQuoL77iFsNSDH45lxNzXcBUoXRKzRsFeoubqPe3Nl9qqJWFx+7
P1QyX0uBDxs3XaeLIPEIm+5vlqouUa55mgDUqKtyIOOsO3Th+DNhcJK3keApt94u
qv7EJrgUPNSbJckiemllyu8fSCg0Ea6h1ImjK/L4dPFnTZeVtbzo2j2Pxpvfs7MS
0Ex+1BAAZlNizuwKExe/Tpb9t6HsYqBSx3VQdFSYVbucFbxeFEeH+Ywij9phCaK2
RD0JwUA27COW2MjQguPzlMJMqWGQB5BqXgXTTrGtroqMmwQ1y21HmH7GFFmHiKgo
JAIRcc5wgPuLOueUMMfBrVf7i73vH0Zaw8/40fPqh5nnW576UUL2yFqPNWwB77BR
gKHxlyds4oDmq7FqJgFHNYqd/pKXbusr1nDhcbG5pCZ0xPY8L3ybYD0yEo/TQqLH
HJoY251xG7Ks47BWyfG7lEj22Z4+GzBWzrl0XrHOe+7DLKAtbo7MbAkU7xHS03si
JR4WEdPvvVAPPMIfDoEJ2t5sn/DJXpj89rMSZs/HRTCRoiunViMRbzsgO7JYVjhE
VtJqI1BPX0LRCcaxEOMhXBQKDKRMrMMid1bmSodMD553bQVHU4NdmD2GYXDpxClh
Eh4h+eFKuLzUqeCvs1NPpDJiD+P/x5KtnkZE4P57a3UuN5sBl+v1zV0dNbiOH0C6
tp69IbyHjPUH+q6BrGpKCVOkXqAhLKedl4k4Aq8BDvxioiL7De5bQLpJZ6l+/BDz
zwSEP9gW9j76bc6MAE9wf56/CJS0roPyKwlPf2ukGNXJJvsmD/oLKM8M1iJOIuyC
9UZTCLJVpuJX/BLZO3371+8SP8CVi6k2OEqICZDxg9KvnAqmVOb3t2kHLSM8F+MD
gVQ3M7c2YKBtH6pbf9COnHLyRpWAVhCPJQhgYjRvTgYDNComtThJNPEL4ZTSsnPp
cWxZCaeaHMz0R/I6EsJM37E1v/EXZnvWRK2eX60tEilH9x1fIsYMiVlaXNPQzrAc
4WEcFBZYPKiG+i0Eg2WU6ltOAHREISo9DJCtTq7IhWt1hd+rL7Za2isevuXXBfUy
fhwUylrm21gSC7TVv1h1VHbMRs22g/0PUbyPKoXxPxHo3bOsOQrz5hGa5gDLAF3T
PtYnverUet9xx7ynYEP93IMhnzB9e5VumsYl5oGGwKlH0cnzzeO79C3v1DEjxq51
S3dr760z+cMY9uyrksHEjfedn0DraBsguvj9OqpXxy7lOoDwunuAKbe1gfHi6ldc
txBiUNsGSv3nN2rLSdSo1Zwzvn9x85Nc9szo5bUaV7J2gShxthzY3hU3gZHFDH8M
y9N+Rl+WCdjx5z2O86nBt0JINpR9koryTSr2XacUsYwnnx9f9pFVH3ps5UlddHfh
9ib2Y07EeFP8oF0k5OZDLJNf6ZP3yHdjg1koKwWjNOi+PvYcit9iTAupeM1LPwMt
G7AykzdHDz3Et9MJyhSacNVoRbzPPjieXBJrFEc3NVwbeAJLvGTWc0Iuq5sw9oX1
ydGQFZpdY3/4/Escsxe35zDL3wLtc1h6KYm7/ZnxIIEdUH5o/aK6+h1uJ03VH4G6
QMsVhsGgNpbvKStxg+es+89dc1Ty+qVNY+yYUgkE8s+9fQoeXIp0jCc1rT+l6xcK
WAKZJ1+xxy3uH7lJTwEN9DZfO+KEifrpPI9Eund3YqCFbVk+YMHj/YqDvdMAfNIx
Np3iIfXuoKjDxQ5itIunwtz1aNFITPGyafDEWxMg/Wt79WmZW/D7AABtOcwuWB8o
95mawtSgg8kNYcmx0+lCVS5cH4KS0KNPKOPe3IpjkDBRyE3ENwBI5ZZFpRfDNyyu
kJmP/NLOuKSkP3To3ZxDQjLt3FHWdUZWEfXbRWAeKiq65J2nEnPmJGF+bsyK4QYd
qavA2pjT3ydKwF36DhfM9kHx2PP4ntk1q6NSbsiPCEXsPJhdVucfxKIUyBVLSBGd
dxmrX9PRNdMtPaTe0SNvX4k3TFkk34T/1Y9+3h8aZFt8u7BXNpmZ7hMIivvlDKGL
mMBjMBBZoa3o+Wj+PG57tlOV46JRukDajTCnV2HODQ7srQD1gqOMpE7tQ1s/RE1S
cavzKyEXdydy6hN2K7tZazMAooQcL3ppsuPFaIX0ei5cQdcd8OqK3JRLUmOMG5i2
0mHxfALHdWq927MFKjrQ4ulemNKaicpT7R9gLYWWVGYSlYt+NWhOfewWrbNmtIB5
/sjmWUhTn3QonZvFkgwbTYDd6EysTIgKvS98pkcN/aBbVSxAmP1gFl7NItpSisg8
GyMqgjsYBhxKCbJFdfPPlQMUYEWz01fRAJrLNlTbvlHptARquBlPcHakPNcblutb
c0bDNpMr+UD8B9qzWwTc9+tX3UQ5Q67tjtP4dBTJtvibpKd9Hz4iCp9X0aCGgV3g
9pF0Eza0w+L0GSt/mNOg3n78yjvhcv/nybTP/lMjdITvQqsY0ng2K3FoNlUD82Lq
of1hG/bADEx/aYiop+UjYTM229j5ClU0wZGnkQpHzJ15vqGqZchaq8XWhLJPieXB
2NDAmObJPFeoUyGuYmCm6H093J3sY+2KJW+TNxXZnM2yt7R/7QpFv20SaUjBhXVR
uubXPFZEucdMZkDh7x30DWjbqSP2Sfvs8oF7vnWk72Yy0aRPDPNX/xMuIQbhwkJm
CI8gMk3yxIUBfsm7hU1nRrAZ9Kj3uCQPzHWtB7IzcovdgwJ3JSSlTUSyg1ZoF2Na
CnTJEIQTfMazOkOlmX7EHoXwT/TS4yXp9EnUzZPhOY1ZtlOr6X9v7fXXuYCqj7tU
Dd5o55oNx/Q0odTralZWb4r+04bA49IKCbFH70erg+vpp2WxRXxAxID+TstLFJ4V
Wzg+eote9jufau3FCsXWZhN3lle4cSMVTqpXaR3aakDVm+EZYygga9g7hJcvSuwq
qBB/uxxEIPLbgnEfBx6ZEKoMytYvcoswADP9Sy41hRhKazXhbQsddP09fwSdrnyy
`pragma protect end_protected
