// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:55 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
fjUHhEdUwhAWrunEiJNVoDa9Kxlb48I076vIfSkAN0dBNiNQJk0CpTuVSemEty9m
hOrf7IqfnUzEx2WPAtU8D/uHILmb72jRBw3K/pDInp1lRC82TdIuDK/tKTwQHbsE
KzxH1QeFwlF5eiZVBCjJZACXyCrmgQwiH7WwRC5vQfQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5216)
YfzPgg10C3VVKaBNVK3g3mIAnywlQKTk+NmD+eR/YibBzYFXpk1Fn/3MJ5AA14ZP
/ZWOUMpS5UMZlzqKSPZh371XH0iMu8E/ZIa1nCdZWh2RgtjOYDriPHukj6ZAxTJI
9AIsMxER8IslnFOCsvAcly7VlC9kx9MDglus/Bct8odxPkO0cuNkn4NR6qlNvNCo
KhUe0rQGLpuVLlL4TzXtSqev+0z4VD0h1NINpd8jDSPQ9CL31/qAqM/14dr6wQy7
D6Tt4ypXceRS4aBpWizRsfnISZ7C5jv6dOwG+IO11jhLwND/8n9ncz7xXNfcG8bY
IoZK63bC3cg1RsP2CNEPCFvbfLBRBQteokGWAyXzsjIrUQ4GKmOpMEGv+gjFUGId
gvaTUtr0bNmICBlF324CRNifSsoaUQ5njG/H94QtDSjo/sTqKFhjJXaoPHGSvaE7
UD3U7bON0Hi0S7mOK0T9R5UayFFrrioDmkNffQD6vRR+6Gl1KQcGYEbJo7uq4DHZ
BH4Y0tEniMajPWxzr2QB0+qKMaB7GdIcWPkeGmoRtpbnZt4jBeZ/MK6uCayi5zbn
1Ee/Qy/9nii9Va27nvLMTJeVybNCbpJArkiTg3RWo/IbJN4aUetrOhB6J64ozTXx
rv5AzPpbzns9uOZJ5nhRbGMS1yF//bjzuyhbgWq5gWqjmaoris4BiqOykZ1RIdV4
1xsWpA6P2aQfwalC+o5k942s1qXCcCAINjYvdu/Godb/qXK3nzYa7p5LOCvAymZs
OqlYd9HH95yxmcyjAXG2GT74D0CWhP55WrIDCpkpIZtYB7iZTeMkyR569IW86ZIC
zpnD0RYzW+d65yVxnFQBJ+eTRlxJnezGiCZIPWjA4N4X1SqP4Qv9tnk/gmWrWHif
ZCkkwaiagiVA1lypTlJyQ2a4I/vcQpJsAWmRddVALoXbX7GwLTtNKQVMPiuTqkNB
jPNOhavVebENL5CYQb61RrP28OYQYkSe9viWa4/r26RIXuOtvpX7QUFgjkkPifB8
vAXl4Qdzz597EJxTyCMIFRtallLIAOc5gMptqxZLDqC6mgVeVG0WCNr8JDb1FXlE
fQq0pf/Ph1kXY2sX1S2OE3Kql5q2szlVrvhnPZBe2nKTCTJaXVC+3/k/IhmmQRWe
uPcVyvdDtoqqMG9bfe886xIs4y+ivF7l59G5i/wJT8oJ65ktFCP/dvZluZEA7jkx
cMUFJ0Nfvdrx3Dqo7ztRuE3ROyjzX5eQfV7wWc9rCJnOtW7BnvB8b+Bx+H1qdnEP
OUZ1LKLMewV+zkIws71mT0cBzAEtmTn4618dOG1rneSgT5ajgLMASL7cjd7fAYjb
Gxc1fClTRvqmGE1zCX5KJQfp2fbuEJOzLJyW3AXwSMkjk8i/ts8crdqW5Pc49L02
mDjw1WkYSlcFAHZIc2YPgb4Jm6HqsdFcZ+bGpasHelKKfIrdCRJBCNNNwgqgYlun
zt6R6AtN2TFOPrmejOMI5sb+3f8Sk7hxWGKSaAZwEOHL+GD7vSWVAnKdHRV1vo+f
u2W5BlJFMwqX0XVqb6zDZzLLjTuavvMANcQzvSiSc5u9Ebxbq0DHbyqsLBNnZuJL
l6xmftaHJs08mO9nhYlaVFIDgOIWwug+t+Jq5BhwU6OXUJdUs4bvv5saQfE14b5D
pY3vgEPuyjyw68g+3NKENhqvyFoEbsRkFjfMFNEphQmu5Oie02ni7d8P4DXFBBTN
sVQ6s2Ri3AJjG6SXnngvJYxdx2JTivpTEg3hPuAQ9GQ6YeQZn7sWdXREddHw43zm
f9BRnKsr4SEZnONNs9tbZ90YNjjMVwTnZF4/9cP2WUscD+DSVH2tsZnA2M6uNlY4
aQFokYefcFpTZeh9ijkA1GR9OX/wJmZwTI+X6XBl+sgePmaCN45rdaeVK2g4eyEI
xJRHP+/Ih0FoJfzfegtGuA76Mb1sQ80wUYEeMVjrorZDa6BgV7qKIxUdjmMc8Cif
texeAPiH/SUV1jU7yIsrWapYfHdSgn5JlbeBOyT8UTWeGk8zwmonsNPKDJIcOPa9
RteW9aSl2u9CirPXBM0yazDVQkW8IbYWLJvqsjYqaibajh3fQZArrMLSHOTgEqNY
BzAv2SvZsdwAZ5V75PYlqbOI4izhSzEjnTcb/92p1eh/RilsGHTgII3d3jmj37MI
LuuBX0DwtUM/Eq3dn9qEH6WHoA/S9g1uRiR7hevcpVaqVL+wWO589MUzwjAZvsa8
IfHqrMNjE8VfoOv0uV3UOhCg033701/D5Zr+uH5XbOV622Vir8b5JqV7hEeAsBy0
Wikt/bC/BlCI1mEpiXwS+I+65/r3LHfiKfIP8LXjtekWEKNbxCYtQ/7yLveaj8m5
SdpnFnM5qcJJ0d13uHxQYgtCQ6USO1eRcvut+aiyYuU1jmcRQ1ipQGz3zu5bguSq
8u9CpD7lTk9Juc+4ooyunWsDU0HZehz9lGwIQ4Orz/3OH12FheU1dAlHpxV/ls73
GpStUKoXUFJ+Fbp5zhJnIrrvjbEmHdQbonfEji5623HFPZ+EADZ5clRRuZ+IYIAD
RdUcg5RTDIhQ2Gtqs5k9o7WX8Dz0SezidqQA3OkZZh5Y/hUS3WzmjNVmpQlky0ey
ZIh0E1XH+vzF3AWBGPMjCkGyPYmAAljDRFY3IM6313Ap+zo1BVtHm6QRA+xy1Y1f
tACW2rM0PBfxUaymapK97aowBpafn9cUO4uW8YsG0LQot6wADcd1OzjXFiw87gBd
hA2hB63q4SmTem+2WfxRAx9OZrcPzmPfJD5t+lwBVwc3ArINdMm9Jtpde7h/m9Mq
JNKKt8i3WpDr5OlF5g2lTf7w0SPJIvVLYBeuUyXFtBYTR3hU3pMvkxvjymwQMfFw
gZeZOibKmfkSS5q6sZmBX1kzI/xYUHOfVCqkDIWVKzlXLe0ZeF4Ex2jml8pqkc4P
PVroWwhAkZGdA0I+FeUe/b0+Xt8oy2yDJlFsciHQJ2JvM8Oli0ayCSytrhTD83o6
0WN7vGGWqDR0uClqbLH/kZTkO9kRT75f9vaOGcEDEa+70Vln+eIjTHc5m/huw9OS
hAwf7ghDIIlJZDtEcMLWYFqshlbamt4W1fUw5XLeBxKRwroLgRlgRo24L6EKNbq/
7wljHvbGn0qSla5OtZIvnY13l1N3mLid/S59Ww5baK0CXKiPulmfOPXEAZEW2Nmv
wZaVNDAnw+PLJOkepQh0U0dVKnponf0sVs3+TD5ea5SvtGI3ae9Wh2LLwiWuGyrB
IbozlPhdEzz8FQVOWkVODO+EhBXsqZUb5LT9mfVQJP9Ekb54jvHMYYwiCnQnNP7m
YlX7WdMvuvX76u9wZUaPF79gAEfrwFNP8pSwOsN7Chx1sTK6tEzbi3SgA5S2Mhox
POI7UsifyPqRsAoqvwHIl1aYm/yffMykUFphV9n/k/Lg4IwAumschpl2nGQ3bkFT
X5uN7TNO/TCAXFmlZssI9ZICstGXSWx+/DzqcfzlLAKbCbbadbFKRTeOKvaGp6WQ
+AQzXOADOOdGgvecSKGY23lVqCLmGSJEHZ1WZbQlaxwdoVJpB1yC/VfWLiyps5fS
d+yQbsU7h2v5KO0ABnSnEMuy1tg3rZreM3k8sLFinlN9jCToqZawW6nmNr3x4378
BoDUDWSnxGk/2XV/uqbk6cViHLpaxbkK1w5OysZ9wo5Xws/CCOU856SZngEUBWpp
meoHyhD9Rfr8j52kQh8O73iM1GrDvj4Mlyf9QYB5wxIkNWLwekvAimg9H3KGPgDC
pxNgzeGEGtyS6ae0T1J3WkXSXtWeGuUReorJ241vHfxXPlPtKpWUnukpby05UzWj
CMzYq3h+QA1yd1M83Oh63kZMmKSEm11u64PI1ew/Fd6yEMgElxIho7cNmkDIv6Gn
frUg9sWpY5GCpymDiMmUL1mOHXmp4Mh8s0pkbo4FxK3wtwBliTSM6zWFZ5I54CAU
kHK5+Tedg/aMLV3tsJeGMWYyjIuu9g94uDZhN3E4i8KS1FnTI4EbP5DbblxFJhIr
eZMG/ywpYHAXIbGTApOYe5mfnKeEsUvqPW4hi5slMCqmJiA43GYMeMSZ6bS2DYfL
eIEjpnJvUswTiKhe/NNxU/tjxdCugoT3q295/a9y/YjBkpoIe4itxI/MV/2o+3FQ
paNvwpjKiGHadOhJcdZwof3QIMfwaN+QpI4CteqB9UVf+vigeX83RTdEwJq2xZWB
E7PaC0ZhRuY3u9XSwQifVC+PdBirVGwrQpa+xNaryszs8YQCwLVc3l1EAwq/J1rQ
p7bMCUz3VMOnIBmz2s4y5OiJc9Q26Fkc37jyF3MY5SXFSY2xxhiufpRCaHJ31sJS
/mlAs+Hd3cmYUU74j9ADuVpS3hsWprdAAOT2QRULPli7KsDbUiXPrA2AaY90SRAn
9Fcxx0LdJfX1EM9BxXXkLbEMZtrKIo2PP+hfFckMzwXzgczNojQwmXLRBhAGDO5g
zsIEsfmOajM2WGJs2NXiHREymwwjbYUe6YdingwGtBnvAJVlh4XFFzYmBH8HTH/Z
4X8UhQwAJiByUVioiUCNLTGk+WWepV99ICXRq09qMTolz5MGjJY6K1mfY+XInKHH
/fcdJGIbJzsHu+KfyJGDwkRyhxv3Ocx33ZYgv+xN4M7oXVSv/3Qte4Jy/tRMwcQk
4sY1vEQ911ANCG81DuKgnBSRnk5f92cTb3tP3qR0Oegocqj5okyM+m/Lo/Toe8jL
S06PEW9cxuJduWAVPsfSm+GQLLHqvuc8drFzEtb7Rh2RwbC9jtbhn5eP3VeLnqm+
c6Rfve/PuKrtGVfWn7MMiVv+ui2gTo/LscXBiAIB9Z0GZnooJXQq4EqjuTKG9KRR
bfPuHdMe32QQz+p2Tc24hQjbpAQOTPRNrP30KFxCyodZ1y0gM521/NV9rOohaNn0
s1M+j0H+uFkQiJaghS3kcOOut3IxSjyrMkzfUifd+DM3kfmCA8YgsNtyDHD6dHPg
3/M5dPvgge6h2z7xrpmC+eUEeWpwq0pwG8wKZHGHR96MMoFcA1ryanoTofwE3I8I
iJY+DwcvVdDJGm9LdLE1M3NZE9wpshWmXZJ5kJ/GqsPeTAXsSHC49hrfR+ZkhUG3
79fYdK9kxKwUrcUQaDIX2tUz8AkJg9ZaBoIKC1EEGt5ItlE6falXXg773P6qNum5
Y3dt8qaXDDlb/hy6K2JQ4QNgwcnJIzKD55imbLnSWNOTGO70NVjK7KvNp8IguxAw
P1cmItl71o6ONu3Tq77jlHuMy4Q7SDafXNQz0Q4w4CnNtG/HnKVItSbXP7Df+Nx2
iSFQSaqACxYW2eO6jUnhIxaJKbybTe0uz8k3F8EDsJ+SrhDeOSLjALP++7BhPTLi
b/lXlke7qP61/Wh4seUqSIPAvnPtoX7fZutPR7VRDoQ4qOnsHTnMS0QD78HUSEuV
QPedcSYAXhHz0awTJilguSeoxpmlZRKfTe+9Fx21a9Bt8mqDqc586maURqPMJPYZ
iHeWH/r+yhVXHsJD6/i8XrsdgPD60gGWXcT0loVqvtYkA8f+zUMbwAvQf3RuDqmn
dWrEcHGQ/7FtrLI7ODlsD6zqccEHL7HEekCnfKaXoXAtQaChGYxCnJ5S9vpB6z7e
ZnmeXKQndStwE8+u/my4LLpzlOEBDKeli0XCTAcllMrpF97+uIQYabakln37qN8u
sXxmP3TZ0TKcsIpDyVsj6Jap9Zba//aULqcHWrULvzfZeJV2PKDXXTCelveEM6yR
yGXfq2yqtzk2UzIuOsPlTF4QqXo/YYguaTUvVnzXHBLylxw5nc9h61USRzN6oi2H
vs55IRizGBEt4keo5TqyOgsfIkG8HHGs6whBde84/06hwNAJmVQO8IHuBlHt2mx0
7AQnnFZ7HiYQx0C1MBUTGUgBiijWjmykZrg8SA+7wBTKZQ6IJn7R0c6wesqR7yUn
htNN47AhYsfyGh2q+DnXPPzbMOIOLbHILmsv/RoopXRPdhVUgCsOl8twE+NaBVK/
SyoytLRaPPA/W9e4R+z1TbjXe2tL0/xZGAFuybi7BQB8Mu3NlnRNcQmofw2+kUbP
rPVT4KmkpRkgcwHwlUDzjopwkWAnrLXrkmwKVBiXn2AqxtV+ARgsp+yV9goqVRqc
u0Fdgoqwg8u8Ugfckr82AOjz6tMHtcNR1KvNXrcgTs5pCYpdI8NxR+HBOiWq+7AH
07L3xOdRb9bInUv8BLkUcKgedMUogaaaQUzQ43GbMCQXoaDMC6wtg37xjSauIf90
2ZxFQVnHehigxvj2+fyqQk741UJ2cfjVMGlkjzJZp4+KxA+/w7yprUYNKPOk11sH
rvP4hGEusfmvjaUfdj8l4aXG+DxBEqcIgB2tm4dJnvtjUGNzHKZSMJSEYPDgSw9z
3JvU4B1+dfOTnnM04ukhuFKfgsobcxDYfKmvB1DDJEvGYPwWp2AKGbpTFUmJEpEl
uAwNFewWZ8blDcIPzRL4nyDRbkVvKjxpgamhwd2W3uDqCpR7bChv0YE1V4oUTUCS
iIgDFuGCuf99rcz/tkYpzIiAjc2sHNU615Hi21DuDET6cOSQhLjX8hHRwu0ThbRW
IJnE3tCBu7cirOYnVlwQ8m1G8dH6q8casYrjvt9RPdron4yA9kH7tFGUcn4H4pTx
bIZxuopnxsMMUTqE6H9NNzyZ4RifrH9RxztbocwlRlyBOJxXufL2nbxDPmec9ekG
6hRhIZn5HvIiPXHDAPHt8b1cp9bJyPFjpeXR05/mCVCOA+YV0SLgkRQhv1pJn7lT
KwxrURvrd/1dRuYewbUQJ3J20dxngBSdTfVtqVFI0wjDVyl8HQgpCYzS42RX02YF
EUuUqLDW0L7PwkOXOZaeBqcghBba7Ae2B3L2oVaSbItnC/PmcSUJ9yBCRsk/Aib9
sY/OI9AXpg/JzGSMN47skmIDAoEyRBdZvXPhHaB6Nw4=
`pragma protect end_protected
