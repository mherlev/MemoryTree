// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
/OaWGZ3E1GSBsvOnsYr4d3QzQ8nWiYiPrDD+Cfm3L5GO9HTK8J+P0JqGe/QcuC7Q
Xn2+RjfMZ5EQi7rrDB9g1fxqSNon13fR52KqablJfCkgfXydxv5BOBXp2v22CfC0
JBWnS63+bH/QcdYGamUZpbqZJDQqwtzYfxmh2os0IARLUHO+JCBm3g==
//pragma protect end_key_block
//pragma protect digest_block
lG9w0uzx5WmxTymtA6jJo3OX1zo=
//pragma protect end_digest_block
//pragma protect data_block
G/DzEF7QzNUuO7DoA30+fGhj/TICA3Q3ujaKHQVeGPcL+wkDYqtsloiItDIC3rVk
WpyYrbAVDD+F7yFH74aPWVQiAIGPuQTcrXkZzUeD2S/pOPOaEvVVyeI05snXZFGG
lOijN5LRTo1NuMtLfVYL94CEdIo7jqY+ra4D71Vjy5Zkkl7pzgjsJlrH0vCJDuf4
Oc1AZT4yBT+neh03zubfeelCef4AfTaplG6c/YqKACp/ap6GeGJrpL//B8fPewxG
CbkYl4JZrjvEK7Y9gGG/etMBRlwzTocfc/EyNzrsYAYuBKpFIPJe83GIM7ulW+Al
YnJ6ebh/ZxpJNhtQr4HM6BzoQ0nhKSl8un1uoAjPb6q/DHuvqAeWtWFU9cAqvAMe
E8ETxo7riQ9xNjxfumBQuzZQ1WMYltAtkJdPZ7VtYTDeq9Jo5GuL9DgeQqj2MCSv
dC3p4WjQPGKV7+2f8Z3iT0IJqGsd8tir7uLe9CXtBTdiiJY1mtPt82JbBAkqkeIL
kXreHFMqKV9UZGnEbCGePyhgQzlSz/068JOic6bbKklbNlpCDgyj5cRMWrYiKI1K
x5+YwQ9BXpOxyQjIhL8Dk4ymlUimWRSF3Hp8GpQpEZhOF27eGO7LQXNFy8yFeiKa
u3LrIbtcWx4Bx8g7sqoIJRcakWrs9sbFIHcm70RJve7Rpu6RCR57/ovekuaOlgTr
6aiZLQDLqlm9oDYgZKoc8YWZ+Av6D7YbTpS8QGOhNxvBB9fKrrZBTF6QmIUygB50
40kAYykzZkf/s4l2EiF99a9VQ6JpjhAMgTeHOqWgzQhfJLzXMYMfdmUbRygjSdfI
v9/42MjzteigFMnKNm56mgy5TCfWH6+9u4/4RTCx9iPeY2dcXVaDsCffKG/wLvit
4n9L6yhu+AwLTDBFfoR0vdo9qpkAFfR/FaW/N1Rr894kjIFAbcqTOWC6iatjo3hc
53T5DMVCdzWapDGiaSfKxts85+falnIEe3X0o5u1S2EzzJm3X+NdCCMKB1Qi7awz
uJnXUUK/Vucd1Pf7hCydh72xOCisZxL9RXD3v7DLGnDiEe9QnbduIP4iCGI1iAkr
W4ez4Dl50YZjxnA6O540khmK+9hP1l+cb1aMw8y3rH1aqhhKM6/FHGACz8/zDWsY
czJFsdQpP+b1XABAqmsylmeCKEh7dnz+qDkYHxuQLXqAXyV2FHR1KxYxDGTWGlgZ
PYyuQcnBZXnzKBFxntxy0b9iAnonLXnSyC24b7u4faCSDRWpcaIMiMZ57Leh/UnQ
evFdtd9iNPalVMuk5uPQ5esmJ0weGy0jaQvAXJxFAtYHbwboeKjnxQp8JOSjsxAZ
lkJgWG0uMtLdSzXAeMHAxVbA5fQ26OuYRU+SzvxQ+gz5Tfb9E+njt8SBNkY6OxVf
JqGjMLv3EpLcf4CNHHb2ceyGnoHw4ohFYm4Zf9mD98qWGn6aDkfak4og8Sc+Ij8Y
x4E8Y9GWtb2t7M8JwHn+c0JO/yiwOYHSQ6ZCau3Zsna9Lyax5pFmifiLvR226SyS
aOyuRRnd/T76rYbqCvaIqpeMPQTrmh4FqJ0kPj7BKBgldWCBCPiwKDvMzTgEaPBw
Z8UAp+2kY6r/GdWAY7EbAD7uHILJ3cPS2RfDaKKKBUYfiY2EvIcpktpXD87FINsb
ZJjtFvnDM3i+aiT/uosKQB+eBUsa1HwkGrhhreFZmatHxtBDdZMwv/9/9q1mTviW
uL6NsoN3HqJkEegFQASlWLMtG8dviJbb8TAIJZOHXqZvTAZszc8tmqs/9QmRhv98
r+M9FIuxescz2WlORZKevkApktY/zSI3ZADHwuwyrH+4USq8W8tbkNXbVF0I78TB
YVQJ8Om0nt1vd+eMtmfnQW/Yr7dNd2W8WU2m1Yg8RQkcvEc+gPeVTWoCj83fxBto
bdl8xVTJuPEeGdORx7AESvlb5sf43LOy4DyOnXX8RuVf55JXs/Sth3PSdSQhllZ7
7OXndcqluN6Ytp65XtpxZ5Onq8BDuq5w0rFni3BCL6SMvvACIiTCI44wtIJtjsR6
f2ElRJoK6aQsrsSjB/aHx9qaKC34uLGpjfgnRjRy6yiS8vJAQZEJ7EzqZ3DVM+Up
rEyNwuVJXH172XEFI+DYP6o6kh7Tt9bFdgDmF9ZUtzfKfCQCqt96MrMmWJrIWmfI
VfKGRAedGLrjrtaGtxEwvEcVcOIEUQtyX05pYu0ERTmYolrUhkd71qi/pXDzIg/r
/fUXa+lfH09vlOqY4ICcbQFJwr3ZBQ0gK//RlPWyEChGdKhbLU3m8t5RE4FYTi33
5/VC2f/oNFlF7rDOGy1H7R4ntX9kRwlLoqScMb3VdDkvV81Ns4LsRWhIrpwNYFnY
slOLoqDoHMTmfg4GT6FGxgm/VhozaDotn5DWzjRpLmlvPOhndrvGcpujl1sQuZOU
DQr7NT44jpl64Yse7b5tF23aJ2wlJIU1oDwUzxXSGeXJ5Xi/TgHTE8zECXWNjBRw
UWN1gyZYEt9RQhwb1fpAq5b4XkpSUdabVZoy7tljrpc8gsrKqpSDTk9FtuRHQ5sR
J0eGfodYI2myspg2eUcLv/NwAAWp0huPowPOTEugEXPWYoq427dM92LyKQInBm/V
rdX6LswYtrUpsFU8loHSBtcuzlx2svquMmvcup33nTj7vOMuOmhY/Bi0bft+Ntlq
Dv4W7vCiSKhnxALO4F7U5ZQjLVDW4CtoUnrIRhYWbRLTf2E1EG3KVTR6VjUurHbz
emCdOoZb11kaNlca9tNcwm1iYqlbJxbmoJJKONgXhxOkgmukM6ICPD3VWW7rB9PX
aMed29Exjt8IRq6Qhfu440K2nXEd/Wwi7Q1IHQzdk6kY3DGAxJDCYOY7zBVSzRkH
Ji/lnowfF+IpntxZT28BOJ4rnJTwSYJ/s9sF/iSELdhSsatfqHZatAR9Xs2UNBBV
ewIm6y0Obn3jPvdhM40FNyDuIgyvIXkpT6mXeo5v7oPkc2UhTTGc9MC3IMDYE0A3
G+WzeGtoRAGGA+NP0Y5TdLTagm0qirz9Vl4kWYBXQmHB+MRJOXUfAqXH99ziKzg8
rWmL1N878j5Sk+zbQWBbyNhdnGplA8Icf4eNjReFnmPks220RExiIADcWBwWg87M
zovOaUn5aiLikN0yVRblti0DxWRmT48iddeSJJGgg2ilsqb0TBY/A1AB2d1/BY+u
yK/aEt/jLtPAIExEXy8nPh/UDXNe92VJhXv/xojULPUJT4VHp9gsYnk0KZuWhey9
IrEE3X7HvCuF9ha3zB8GmJ1zYU+09AwTs1M0j8ha9n3M3PFOmeMTem+xw0MMsJyU
zuszyiAWRq0Sx/sy2y7QPI+wnP1JrxN3VaXj7OKBJzcMxddkrXNlIV3ixCaN+0mL
IkqgeF+s+i8Dgm0+jh8wSAwPnkOhYnmQrjmgmfIUHytA2tX8eF0B+LgjJ1jX0aaZ
IjshQNKabe0kLMo3pIkuXF5a3R4b/6uRQBSdcf8iQBQLN+UQdp/p5hP3SQ7ju4ge
GhYCXPxuBURnAxe0dSxNpFykyRmq8TLQI0fEeWU5LNL9nvB0X1qGYrN+ok+MAv1F
R3yS/6n+9inqzP8gOt53labNlXW14Z9SZz6NEmMoY23dhcixdMGbcjss1/pgQC/U
yYAOGoRa0TntJHrE9rYojBxokriSmQ+u5mnyXmUZOsUScuV27TeAENnQ/LvFfY5X
sUaPMQZc9z/ARYjYFvEYfF70l7yyPUFf4YsMwRtN2CmK+ZgnWXJkg/gvhYUOFZCS
+ylHRGEF4ES77ubgdlldf888iINWK75FcLmQYPGEY2OgFB5YooZzqkEH9Jx2Tjns
tD/AjYDdOSbiFshKMC+9sZNEbaEQdLvNWu1o5hDo3Q+l5higLyvsQa3xPoUyMEMI
YPhjWegUnn6tDf1Go5UFkT+tsjKnRIAAok34Ggiyqle79xNE7Sb7qw+tBxoyssB8
WivN+9ePb+GqRIEwiGRfa3IDDI3WFG/iRTVbQvEVqIO8g0jfEPtghHF2iDEpP/LN
dshUKxbe+DMW9pgMPLsAbGTImWQzLnkK7+eEwfXtw0kbfXNrrYDmCCpcf/fug0Jj
U+d2Kxz90SBa4lnrOrj22RMrLvm9+oYGHxq5HPsr7kys3QYwMZAr8vvcZxVJQ5i/
8/U2qA3X3i1FwP37SjfnWlpTBkXTFaeGOM8aSyY646FeaxN2/2EKuCV03Va6wYzr
+QBrnjjvKwK31V8pR18EtD0dVWbe4Ihtrza6Vc8JYuSR/mm6CA+rcn2gG/gx5kGR
g7eyjQZmGHQm7vo4ehJRjGYS9zZUQ4G/hAK8wqNREgnZ4GVxwL0n4yubPYMcJ/Ok
RxMYrZl7EHXqPyJ5IGBNoxo6r9+RfO2YXZm8R3FfnFaz22k0iYtwRJqIC/s70XpO
uElSRcWNTuWXTj4OQr4Wxk8lXpGL4onVypgKxa5F118YEqaEC3fdDjqFVQEuzqfs
SPORd5stu31MueI39fsKGP3h3DFolUVHSQ1sErfafnCxjcpFy+h9Kwgdt7FcS/Jm
B7y3X+iPxdNi+8f9ii3po/mzz7l2FA3kNdz9eN5uj1aN+Pn3Szsktu/MYTb76y9E
iGPQfNiDY/NJvO6BvGNclqhuay1KlyTSfV6Zsp80BY+sh3f3v5JsBQkd5acnQYw1
rpQkwPgmFqRV1HOZnERQn5VY1+S+xFqPiJVItVjidQwuW3I0xPWf5zp5jRB5DCaK
haPIYtqvCznqSO3dHDl0Pwns8FcXTynBk8Ejd0orZS/BhdXflI3eyZeMaPyBIDK1
wOZ3cK18boX9yYV2F2QaDBQakfq+YNtvP/Z8jG2qHB3/77xII7mFbtbXVVxEiizq
46Jk+UmveM3SXeEmzZyHvqH7Qn9Nv36UfunqBvauAttPCdba13DvY38HGerv/uMC
RsUeMEvlsHlGONs3djFac4sPzct8y+1OJ1IwGDFUYGtLvuSqfJwJ2anYYFUoc650
9P0XhMU9PpKtwSe6jFo9xcGcO3+iP9jPXQhI2CZKf0QBTFFQafArBzdei7ze2qd+
+xF5acwiRJ7HADGC+fVEouy18zAFgvj2Frsw94XpPfmeIyJq1YM415/qwSNJ2AY+
ZP0hK/1RgYePxup1zKIvE6MAkdKMZzPkTX5axDyW3KFhbsVXMlO3BhNjCt/ORORt
DlYAOEqvM6R2hf1iPBmduw/M63/TDgfZ7neyelI9ND/kp+abHj+6PvU9NC+wwZQm
jNxquAt5phrlIMHu5y4M5xJPtZgXNswhQWbgnq+oUTQzKSStZxmzcZHVlV9hfte6
4Fg5ykey9q6QYIabXmEaNdnXO8vqNZgXupvHs0IzfpiTGgKMHMSNcem6RbsNHf0s
BcycFuvKWFjOAgAn5c5844Ap93F8gqix9D6SbyKFjkx9krsmB8P3q6LMvGGmV7qR
fWRxZnyLkt++6AjrvhDEEpMdUTt4LJQP1g0OZsSaJe3xgydTWaTs49ImNmRos9Sz
7y3om/V6o7HD1vvEqYwV/V8jedf7ec3aNjDQLXck4fDuIZ9TUB02hVyM2q0/A3WO
kPSf6VrYikakrno5gqEYGs/GT1BZIN+Ap5RmvOe6hpEINujO8+xibDaecpSXlkDn
4E6+Uf6clIaA6p1AEMNt75Ik+POEch4YCqrtGYCHRHlYX+9LWwkOs13CszJiXouB
Vmr+Qs3UHguf2h0DzppP7mUwt7B9PegO/8+/0D9A4DqNGRWpDM02BExl+s8xeyvF
ZTa+Em2plpAyGs0y+Nnln9VZRV5SwNga7Dj429HMXj88xvgumgN4QWKGMA6qW+Li
5o45AEH/C97DUZK1thiH+eyWaGqZAMnsRT9LNDo+aNsb/HjjYAQaEedVCcWNa7Cp
QPtClCqwChHQTeDN2D0b0M6UT4+G5BRZCwvNS0eUajquOmdxS4Gy8GzVKZuco9zK
/THNv4P/cMSTH6R+hHQA66lXX+d8f3eroJwlqsAPpWsWqg1Xa9gNCBgvlOOYCqAU
Gur8AQfpEMzlv5zl+KqldtlcwisFPMjRtyl1ao+kFIATf4ISYSu6sJ/YZXsH0zHF
kLOdIIq41n8O+5ebxF2kJvNqA9/hSE1DXC7PDJ/W3ri4mQ3bSf96koUWevyKL3jK
BBE3D/tXNYImD7KxS6nCg0tt+2vkATC2jWnId8jcQCkKvcqDJ2P1VV+gjra+SFV2
MMbA+DvRlsU5oFs9E2l4IjPik402tPGpeeAHAQSa80PcN7/gxVRPwi5wV8wrDlAz
ZkP1mBTIPezEgZ465C4utomJmNFMAsbsZ4M5HdQttiw7C8beM9w3/TNnyzikHk/Z
XA64wBH9T1clJQLclLBfGJvkWwYaMkX4Vvp5Ib3VH61xYaArEtJ/G5RT4vu35Kz4
Fm+b8B6xvg68G6ys1hyAIcsSnmL/VJER+fGH0W2a01uAC+wnKHZxUsOTJC2aGMo/
yjvrZmJ+ij9By1h8/hIAZBu+tK8jTEhTY4OXw4XyxfglDUL6SRwfG3U6vAiEaolB
BXzCs0VLea5pNpO2gN22i4uYMSYhQMRpdM15WpESK40iLilSzPOWubO0YjuwbEmf
s5Kcsa4FK2tYcii3vYV0l2ryLtiol8UigUxPtfm+odPl4QxAzStmhcRD9k8BHfHz
Ij/axwHxreDV7IZISOMlDUSXLCFhIOznCee5E+afvGOgHAKdxh8GDYDRMRE/01dm
Y+HGDhr5PWZjr49JJ8svp/dc+fq2c6L9vp6RszIinnGjf3ErAH/T0b4aVXjHVn+b
wipwzD2GzmYhtJTCjni15aV2ufeRpESoMoYJhoC8bSKQBGswc+QGLa0SLS3XglXs
0n3+8ddosVh9EnLUVDnlmYZjnp8mT1mPjuHUF428idX3rkTfNv9lLS34PKRpbMB0
D35zJ9TcFjW+smhoy1fdxLjfZcHYjEbbPSzOUfDovI7zI3vL/PJqfRRHhq9upStL
hFOgzvU4n3dsTQh771zFWPwmjGEC36TDOGF3h6WIu6u6EyNgaw0lIAYO6gaHUkMd
aXfBVuYdibLR+qvnQahBNVf41WTmgaK/R8TmmeeR0DdQsP1cWNgokzHN21TbCakK
YO0dE/I+FLMoCqJIsvFFZTTilkMDnmoYFurFRObvHDFzyEZkrztQYEz0f47b5mQB
vr+Kt6hsMvvgqF93687soQ+/GjRheORyg9uz85EzrklGJgRrhf+R+L166sBbFbaR
XSEjxgrfYurg7rVbT+7uhEValFlCA6kvAeoCJ0w86RMcaASAd+bbMuv3jbG5ZLrm
R32uZ7ISAhOiv54hnXUnq81fiIrb080GUdXJ8IGlOSoqydFXRnPujDLqKeqjMsEn
IdX0SR4vjnLB4mIkQCcw+HCk5BAG2Ap1lOu6eKYf4cT6D2IcZmku2MqYgx4QWuCG
VIC0sixkCfCEG6KZRZEp7UBTZMxfn7TKIua3LFJ5tSmR/kDr+aOQdAVhRoNIAFM2
PTm+MqUX6QGkKZJt+CD8djlSHGOP9233D6KzRs4IPOIT0hnBdSCRfPa67Pxy3HVl
clFPSq4oCp06G+WQUfZV6WZFrCWUUnMTp+f5lKAe1q3fYu5L3NYPBWlaSULrIyXj
AgWc9CqobSVfDk+cQDVue/TmOAHhEl0mJb2PklbxmAS1ew/+PdfyxbVxRCCoZLOE
ieT6TTuAZ34SJo379cIhjRdxKAF5MLyklKEgIdbWQsAhzmyGrXMENEy848TjSLmG
DprmMc3G8HJAE24q1k8a8WX1SqGEIy2YRI+rsG18EOnJbfIyCtYtRYXF8HUnsdqw
bmAifra+bms60uY1LUIgrYGZUc44s6PnrAjMHJveSSwPjhSpDJiyra3jB9JThdws
mf/5rMPf9toJn7IwgRpjBHzPj1UrsEqbOnb5JWKWRAiSkSF91TX1DM8hTZ7vjBXo
ERDPFrmNa97fT4PfC3Oz6HvBGAnEDSYKy9WpAohRXsjzvShLGpoPTwqRbU2d7zpb
LMYbq9qhFCds3vGEBAOYeSKMaLu/iAv2NqFpNxsqxtdLEEliK2aIh9yhsDt7yjdN
Q/M4Hy6CoSwTaAbK5TGoGviO58cdVKVpq+XH2TLzZMer6LgumBwGdKfjbT05BoxX
VDd+liMvDFIxQ84EYlX5+PHAglC+r3rzAHJBH9wg0VjpOp4nYlrrelc2QnQxfhAl
olWGXDIKpfuwv1HCJKCMoghAu01Ql6eBgGFfd5JBAFoIR+MSQ33Gap+qFsVa5mnM
TIgJhQGDnud9KYNJ+pfe3zOOvEEbr0Ye3vQVc8L+dDsg6BFGNUT1go0cEqKn4Voq
g26CR+C8Br0eTisELqfSeDyaD7dxrfgcp5blTM2jE4yQjDlfWdGGDL1vOAugmvVu
jZ/08h7+aiyGQaaJAlJP1pI7ZLUJWr+xmZMM8StbO2572K3ehpSgOyg+UGG3BHuj
TcieJlkypW+7gIUFi1REImn2jP5V0mH4mzX+ZADMmQrQfRUB/sSnC+M6dX/yU1U5
DFUpynYrN/40TJqbpNII2MF3/6TlHwJlZN7SbYk7XoHjbWL/X/465ouvPabFb/nP
3e7/NGHWjCUdwpyPcfFHcNwKwPlDlbNTwnce/GAhkCNrJH9bzuL7qXl0NSuiYtmC
lP6u80Y84lbzrTAmmMSLXYgnC3H7Ds8kJo5N9wpaKjK2/+QLXwgeyBx/nB00mvV6
6I4vp+/JsX8pZLXNYIIvTO3FePJxR+REFjVjzWeQ8YzvHqSAE6Z56pbl3Ah7lRa5
0e/VeSHhFU3/HBgLU2WT4HiIEs0VGxBWmLmr50U50rxDLCl73AL7ow0VEqlPa5Uo
OE3+mbBEggnmj3pHdiRTdeM5lKhJAF9TrtlIqgMfOl0SpNjpOnHAojUnzsbASAUR
07Xc7y9mQOVhKaLltYAoWGmWTTfhtqAc5pj+5SYiUC3+food2vbHgEF9xev5Bnt4
vGKK/cGwl7akAt4k09/v77kCuwWQ3MFO2PfjRH4pCLqDanZJtVRHQbvp4eRrXuTK
7uQUl25IWaTiJgrclrhNX7Tx/r8xGXWviv/rf9xqsdsXYe+cmsYSRK8Y1cgevZ7o
EKDuqglHKjXs9+zC7oUGsCm2Cn1gPPOrfy0NAcPkXZMBBelrPfrXENzWZBDBFF55
M4r8w52INoy45K0vHB1KGyDT12msqvlg1H/Vqs0I4xXw2c71MfWvWopaC8iC3OAS
CP/MczgHefYjot+uAQKkgOB0i19S/XLqtoYKJDsToK4TGvh8D79SPl8vyzlYN5IL
1Wwtfzs2AUYMq+eh6TMTSyH3Ktzi29deSs6xMJKy7VJQ/BiJzJ1bNYnFxd5viY8c
dOEwbCGuLxmkG7TubDoKtxLamC9VN95q7hgXRL1lIH5lWp1qVJUe4k+dJFb1E/3X
sTLlkurojACuj2DnSFha85sXhuOa5m/O0wXDcsimZaKXBoZh/vLrYU1xBuM1CLzl
9h8tIpJA8McHH23R4Bbtqc8EvYH9TQjYhhSCK+szV978royJ574Rnxt91OrDnxcO
keUpppYJAx7Xz9+rodfw0llW1x+k8JFQ99BuuIh8RQgiK806qCKe7t3pQDvmL1ui
Tn//Zi+d9VLWdLwew82ualRCPbFGUHvoCxDu1GrquP2hmNHZ3h000XVCLTjTG/Cl
5HuVQFQS7jTGvTr6a/IdESsMXP2t2FcnAQSlJKSDG2QVmQSqPrhj8D8NIc36BgVo
6TF20bOT7zJ0P8HAZKDWnnK8UMKLWx+I0xbqr+Ow5T7h63QbpkSoGJflmD0DS0gZ
Kt8VoLNPc0vwNRFdmFXvZ0xH6kG6+JLXcOagdWc6iqPHZDTpwkjGNCpN6JQycWLw
pKWB73xbz9Kdtxde6KOUvr11DyXdKTb2jgkit1b/Jis7aTt9F6LBCGtRjTFZNaUQ
S9OWcPNHJpXj1elu0SQWwpLhgBwxuOUfomCxsbSip00IAEGc9FXk6/2Y0IzkF4IV
IadYOJuj+kl/FNoottbMU054SEi8GyrgR1druV9Rg0EprMjRY9xu2nq4p1YGAyRq
f7fZ+F239tJMrwIRygEXp18/mhL44UPG0JmE+xLQDLWlTttHj4GXr5x3WmiL3vb0
+u5UDNezzJ8dw3zED3KcB9cJiyMDNuEZQcFX0ITjmOtxGP/4YJXNAHm5kpGhDzjV
ew8Dee6uarHqv4mp6CfvEV6y0xnRzAP14hRXJdQAZhpcyPutJhp1CJs5Du29YSPd
eq5s7Z4O44UcpX8ZwIvfLYz/vzOAFGzzrdrvuHCPZ8RkYP6rWKOMkQFV8zLwAZN4
WteWIaI0BiOlmAMN+179BsC0PP9EFGJ/H6HTVkvn9ZlTl70j/dtVNKA0fkQcrcPh
eY3Qk18iBN1j2heOd/EWzs2r5043W5cleGStZeq9w20Tc+Atos65QyKXvH9MGbGk
ueBuaXghaqANQDZGRtR6haMJTfcNVTWmhofWdgWAfCxWiHaz8m1KMXlbBwr7s8rR
PiCAxES+MA1Yx4epTj6cFLCjprvQVQXrBjToM8yi8anF2VIvpsUFKUOowhK+6xsO
Ct0KUkYwd6zu4K1FUyJ47+fsIzyqV/t35pWj988HU0WiZw/ktaNvK8mnyR4TZ3NA
1qcYRrbzcpYxdm1QknUPXk0QtHkNXJlLQj3WKN8MQTY47vb4vZhXHWY09mZ6hy6g
qzLJdcyWXYIaItR54c7r35WHdwC48QRlfbuT8KjSiusbnTEJjPpgUcVZLktxDVDo
DaN7Sxi1ti/CkJwsqSNH/PVDb62K24TkiPs+gR5QF+VB+qsWdoPI/AzOwb9LIoHt
+TLfCcgGaTfViaisEPPwkve8WgERdEQS7KmXNv0TqSh9CjU7LpJc5Y6QfDULAAca
/mZYFdP3c3z4ZihG6TvItckK6HF1X45xT2TQA7uKMkzS1F8gcA719lbd84qqLxk0
eCOrtzwz9KNLCp49dpzPJKzAeYBNPajR6IJTYFwIbdTUuzxWeOLwjQEkToiSQixr
XR0ZrvGzIA7PlICno9HY/9usiNOQm+dFoYGRkPwdx7QHUp4XQjhm4tDNFz7X5RID
U+Yqojz068mi3EVRWVAUQ7tI2mQeK63UWq+G2AT/kK7JF3WNAmlJPVvQUqFake4B
gnd+8DftSCB3+6AawY70TCt8bKu7y7ehaAZVRXt322KIBMK96hZ0iz9dPjlxTbG2
T7SBuHl6pp+4Dl4LFEJwP1CdKwyDTYxTzirUaBONvFyp4U55im876izxhjsyXPrz
2o7UWh2r5tdweCxxRuGDYCdzSk6KVkLx6FmC5q/lIo2uLHryVnx3P86aByTnVXkL
q+4Kt2PU861AlU/6b5QowkpRWdc9cOmE5TCZ4VxTiMHWVeB3+suAtmeH0itoAizE
xEvj9GNrgiYI8TsWEgpGfO6ywHhph9xnzZjjhqyQyWYcUgTT3KJgTHUUkbxDG9h4
t4Oi0XdQs/f8/UZjmeqVNstMi76745doBcXTTqHDpZvZb2WPoW/WzZvupiKRi5bG
c8dUs1uIh8d31Phx0DCGFof9hQZqTBcU/TR09/wqIrr+yL3cGRi1I5oEhprrCsrN
ub81irzFELVgTOA3uVHz582dxOv1kVTZrcKYVOQxgGX1ZqGXf1vFnuR03p5fGQGy
QGwUYQw8zSntiEKR9DgNgaXrYT1ZURw18bcgpvfSm8vmzehxdmd7nEWB2r4FpMe7
D4dZLiUOcxPjHUVO7jbHEhHIm12lkZtKEo+U3l0Fm8LblUFv5NODZ1ZKHytRSZej
Cen6TjrsC3y5hx4Zrm5f16s/w2fTWcg0nD4xgBTPLohwTR/CPdkD+yIjeoBbwl3j
Mt3X4RL8asRdoNgBLO9OJf5dwmgoXYM//NvTNUaFSARhuHIRtFbIC/4dBeWlD8MC
+HgbcWBh0X22XZwKfoo1CV6jtGlYloVwMm2n9TF6Asrl6TTuTjMUzSa6n1300tBd
LPgDmE1e/tHKGaFRinvqmHNtDcCbChGTckP4BimKkM46m+BL/6dqo5bxr4LFQL8+
jOLjycGCSBaMrMpbWz2jXLvNjQ+WQetA/Y9LbDHUvXMjqACqU7ImeCKPNBLEqkk2
dqcLxEFSbgHhGPBXUK/AIXmdYzHtFpwtizXBOXNxy0yCxXqjYr6x5owB3h2OggYw
T1edmFqXcSzIxdZnW5fbAmAMYKKuGm3mOkyElKk/V8KFd6HrmBtydnAAN4UWgxN7
imA/Nk0CSmKLcY6UuVodniPM0hE6qnbk0S5wV3eoTir1dDJEcVMLClz/Onj6kzWn
9/hISCYkSIo3+whVxaSsPl05PEg7ErzItMNTX64zehJKqda0Lgu6vbnUQE9MrkgN
aeJDOIDcMqcRUMZnHRwHDV1JwQlVvIOkTXHoPQCbVnocsWFwzj6EYAcutQA/0ldP
O0sxCuqO3mt0KihczoS/DoXB9BqIm6ldftRM3dsyi0hr4HtejQTEKTDD95UPpcqn
C6B6J8N211xv+roWOkqPV3abX1TYXyjk570xkJvcxoX9yc5oVf4DGyHwpOal+BRR
svfpAzGkmVOkjTnspGQyGOCzuerZQhyV4fgRo1ob1+7rJO7CkQGngu7Y3MgLKHcp
IFHZmk6CU4Gr2o+hw+g0V66O5JcRmgrlR5yGGBSYI9X2OpLl1sN14di/1oBep1Tu
xlmYE+C9OLJ5OfL+s9bd98wXlT0NjnhyvJkKe9Hnt6c9hKCbexablm3uy7wN0Vna
EWerW5hmv9vC2fOntRRag+z0bxJaVAK18w9Ny1Xuf3D2fF2PdiJbcdnyStUOxLTa
IEBKWL3dy6X+qekHYvjXk9/S07NK+l0HEtcgw1/NSwF7qULJdjIztv1cEE/jWYWE
TrRe3AeJT3j6qf717KdG9dzuNaVNMT7xqeu2H+7J/3sSlsbk7GXIMsVwHFZZYPSV
ZCjG1yWDwNSII074cryY/AHy7vVB69S94H8u4RqrIazSYuPw69dwZEpRZRTBKLYk
MU+t66Fa+y8+hPfcizTWJ1x8EnsumJ/iRrAlT7vz8yDCYlGGMnsZE4HwJn3wgT9h
ilHcfbx+gkVbR0q9SLjrWuX/VAtHSAjCB0+/979cTUjknmIOmfVWwCY+nU+l1aVp
Z4Y1RwPR21f8HuZsSM5teR9T/1b6+H1GGAABHTKQWmoCSj5U4b/VgOHQyb2Sqxxx
biLLCX/KCMe6RgC8SQf6oPSg+T/NCiQC554F81zvCfspKUc5RKVhgBKj+Rez/XfT
bassefwLj8PO6q0d8tq2ca+0LHHF0MwlUTRljGB7PHlsQ7/3Bqh5sG42gvOE0hzQ
R5kGWBjZvfHFHF7WHG4cHbm+C9fTOuNgPuw0LXgjQx1SLlLV4mc+C88Pi1zeSQzh
0SHgrmGf6R7clYXkl9the3Oe4Jkb5XNlYhBl9n3UewdBHJeD3yBKYn0fio1G9k7w
eqo/PTjOwR8eURey1LVk817RiYMplgmt4vk7O+Ha5MaSkFfSKLvTmTvwB4cY5cmX
lcNbkvlx77Zef7rBiGjcBvfuvysgKmF7capMczbF0jLkXXhGPcIAanoFljSDFnsD
g8FHj3mOoURWjFVMCJYspSJ+zVgcr8qBAs4mAtQ4uY82x3eBIP+pJkCVE/GbigjD
aOBtUMgODwRcZ5bAP8ew2LMoJXB0tgVrOLTfRq9f48tSoL0QKpa8JVJGTRp+18t8
C1n9tf1aSqRhDTxOYAyKvOC3R8etqMkrtoFirbm4zdaKemjvER+32Fbz/07YadSP
sbxHFDB2JMyIbbWJK395K7oh1XF61qMmQFQw2dZdSZNCXq51zUAAYXYjxSQ5X0ab
opdZt2DCmbHrNimMv0UrqyLrxDPBeB3y4n0A1EjSkt1JsoCaGHftWFv7x5fa16zz
JMWra4y8xfseY6gOW+nXa9i1TqqpOhLGShF8g8VTNUYeru6O2UQPXjxXDf0I1ZH6
fFgCXaoKv9Ob1fS+mtUFz3xz8PesX9BmxHJbUpsm519FjeG0WP6pqaeKsbdWm7Wu
GNmB0Agc8VL9yrnbK1cXQOIW7KkzJJs4jQEo69/VrB7Jyw2P/ymgdW2qun9cxw67
JZGbinFh2dEODJuQ23nYvnThEb8BK9tIGjsjE7jVwf3CMIPmEa1YrCWBgP2OlkHY
BArfDJMqRTkXomtNYN1EJVVtNiGQGT0WGNaolTkvygDIoZc+rXeYUwIJP+z+Tyvf
ewgbCLbWRuGljO8yDDcNe7neFF4ubDsGmdYPrbRXaNMe5okWgW9suE6xS7PH+Pzo
DyvGlfUAl9cOLU5Rdr0Imt9okXz4ZrvpjnEZgm47qHyQXR8Zx6u2DbFDTTErs30h
UnAyU/VT4WCyig7nbPiQofblJ2/d6Gu4XoO7WLg4YKotsY4iwRGnxN5G/d1WOZgp
KwhTvOvOx7hbZrKbO6C1m/heIZkASD+9gQ8uD6EaYgRVJlntGxLuXQPDlBfOtaS1
QCfCg3NM+WDxGS0nUrLydna9G+kyAR0f+d1ZhxKDi8Ot0hO2UbCn47cNT5BvgFfO
8ArZc0HhVzMrHOY1dkG+miXHsDG6l0Tf4KYGFbojB6Or1gqY/98UeTxrH/RePWfT
PT5SlTdaPrWT2/CcTtzNZe2nUEw1u9/I9gjFxxUNoMdLfM8IVEXor4xoJhD3A6iX
rbIUxKE7jLhuo3sr+CKQOkqRPK5tUuA8TwEXSEQiBUcli2vq6FKsu5FyjHmkJ//6
WtR7+MceY0mJsOVzBzEm/QDUmgYIO9G+5mSnCmuIphgOVM/kgTAUeoE98PqoaAdg
Y2roYB/J2BnbHrbnJhYWu1Vu5eu4HhkPc5J9pmVyvvtNiVW6r0pPYg0OULunKqx3
/lUGpAl8iCK5FMdshTFvYu8IS+YNSKRnJC32Fc8pr1RVFH+24Kk7UpcxC4v5K5FH
lfiNxn8j+RxBVunbRocMa6of/9wlaJrPQm2VtHWd9f+Uphhpqfqg/v5sxkNWJ2NP
ETfwvd/TfP97CuRo6jewqTgdAbelx260Hf5SeMLrZeBV2DSVpR3G1IWAlMMJ+rm4
8VRIluXUgQOkK8hRZSQkpo7qOFMEtEaAUO6MBW7PBSSiQSWNbwhlT1M9eA2NqDMq
3s2zp3inS5b76x79bxCalr0BobFGFKx7WPa1kIzU1Tk7ICedDQpeNtox97jjE39L
ZY166SpXXO3mDnRNOE5aw05b9hJm66Zfv8Sn/+uiXo/IY/tl4H5BvWZK/b5NWnpn
4uNSpGfzPGnvis4STguIn9W/iImh8YhkvNsbJARKFoya9LcK3ep6GsOt+YRWtvnC
jEc//bQhtHhXi4oNn/zuW4tY3mSrArQr8X8a6VraTARakCkGLiyXuZrRs9vgduuL
l1VoOh2BB8Dei6OlxNSLkllcgIlN1M4jv8cYC+M0wwr2U3nmi9mo89hzUQ9jWFm5
vtp8h/9482yvzQ7N6xQ6qHpBQBv4A8q0RXUcrzXQ7uxpoqjrVOTsklfNHKgGjBZs
d5jTVJ8nYafUGKYZGYb11/qH99YpFeMBAGgfFn13QdtB+1EC51nwHoAHS4QFRSYg
CIVJ/mSdojRRFXg1RcK1RlnuGLD44BrGvw/cP8OMFX9dpz7FNhPMqCptSdDDymHj
bNg4TUtismu2AqG4XeZ9XgjeWUdF0kUu/883yY/APs2VY28ryLOi4fkm5nBsIuh1
REBa7HgbrzOy9k2GUjiZ2Gd1yXC+p853VnLZu1AUpA71Oz7FhB1tpNKGgN5cuASs
+RWdZtFxJuVQgftBQtI8CqzuHPSNoRWckb8wniHfrF3KIPui9w2dsYzwhyS3Ogox
lJ5KLJj9PB4+jGCVlaha7A/KYBkzisSYcZOOfsUoG49uRgMb8lUDKDLHWNQtDYYT
uoSGoZYnGChkFabVCh/n3NydO+NVESJQ0OzhRHZ9bULQFKowUKWwW2/J33p7VrX5
Fo79Ds+Yxi9R6IVLY4F4mU9lyVDbcGaixr8WyU/wpWuypvZn32vD2HBUXar/l6fL
Im23aYz5IbA/SIEyP1vRKZuie0kNVaCg5117O7ZCg5Jt6k1Ms9qx4wchCXI2O8Gl
Pq7eu3nm25mN6PPKx/YDkr6y4M+OaRkug4EmXljWqT+ciijdYZQ5LHbVqzc6OmCl
RHJmQ51H83eWz7u7uW8DRRRz0ImjFfABza9s9x+qAAtm3T2xfWBHBvdu4wv8xxCz
DW4Rv0z53nW388jcB5iUPngW6ILP5G+aYNOctg74H2rmub5i8MZSgHrqspe0RYdq
mvrqoCnTOTkrhSiU0dk+KMFtUI5kb1+Usqb79WaeW2EBCwxSg+l8I63uHP/bG9CD
lyXChO39xY2xc5UYx2jm1fKwgjqQNHB09NzGCA0WLlcvamPjIsDeasALZ0uh5tA8
VoYDiCVWr5rDINJmfpR1iOGOft1/Jj5ZFEG+ziOFijNrWYstgsvCgjyubpQHsJnj
P71ZHT9UBUHe0NFsGaIeyCpRQWGSLwKCKxeEv1/LJofCXRaTMjOmTWcb/uhfK7QD
RT/ANZrYfsDUPgmb560MygGT49mlKaMzN8KVjR04q9IFRNwIIxv3HAlpDKIOplXT
1fG75KUS47B/NMlM0uoBPiGd6j+9/lXX0qMSw48RTFi8bu2KJdbXrNWT5c3Ly8XQ
3+jZXElkh9713AWfH/4oV6exvU7mSMXppCkpscbacvGVUJMyfoN1mPMwZJZemNfj
Z/hVYe5CBZSQhHDP1W24B4DZlhvLn1lDUvINnCIhc5YhcKCq8kPAtWim90HuBane
uomWh2MwWsHU43lYPl62NeMU28g+SHH4XZB+Cie7H2FXzus5TqDRcCK9RK0YK1A7
Aik6hufsS0EpU6XtGhBCboO5nNFueSV6P2eVcQpE+3TmoLGYMYJnOuOKeegVKV1F
4eIIf1HiiyvqYCuty8mFEmCnSRIIskdE9Oz3mssIMwjik79PAPdEGzS7or06YGGm
iGWUo6sFtHlSd4+f7ZXH2f4MO3/X/N9wao1KcmmMk2NH+z6q5142Kg5P1EoErof4
EjtApOaPe6c/BaOzCOuue0T8R9CiqfZhRH/Cpl69igx3xpikEdmTYISYzf4CvtRt
98Piqgws2BgXK8pT0lTwYSQ6S+3qUwngVZ4WZKHXONaVY+YcMi4+qbL95WbP663I
h+XhTlKxR/2Gs23VI4MUwHlJY4dVOZeu7faDknqFJydxM1FO6o/2WD3dIgAt3SBV
T9LpzOGPnKMBod+BqTyCs8NG2+rjbj77tIBqG5KT+QObRtdcWAiuBZ0ems/AdQ07
WjWcTxg54EZFjdR06wmvzpr+00dKQbOO2Zya8QlYWOQEszfoXq+lpEH3A3gFxiEV
R8m8VaLGXr4IGMkmmgJAWHVhQBSR10wdQtLC0Oexun6S0J7Q2uwkXKPnnyTsCWLR
0F99yAhR72ththlTzowBTXhEciLhK/AU6e3zrA2EtFYVNg46AtJ6G1JwuyvYMWs1
Q1VidyYn2Hcf4r+o3ByWwHjfiKkynLKeQdBSs/I3ILNTPRZmEenzJSyiIrrDfprP
b9ND9eSv7zpfije6wP0ZIalO4yKMqEiZtlOk1UqLO60nRI0RAMv8b1ECf8AFnFK0
sTH06UWpploWijoa2vvV6BArZT/egrel5RkKmVSvq7kjGuHDPHrX5mU+AWzmOTkL
UxHhmZRFoUg38xJpjREE1zm3E/QJ4iqd/EjbUUmjQxyX0K5/n2AUXNBq9lIuKeIs
y+FGbgnqoTgCLVir/dMZRwAh4eKz+ETtcASkHEM/4p+yk7KeMU7DqknPTFH8qIdU
2T8XL3v8eshf3Z/xukv7aPofRVBiQO7PjB9gCkVaO6pYyYICxrsHGFuEHQVgJBDF
MaNuf6wZbZW8jLLsoGsmeCQ0HEZLELhIyZGTHKL84xN6q3iY6GkP5WYOqKYnqtnH
u82aABFQpWJmZpo9JtE2jGkNsPRH/AC+xEDYlV+kgS2vYxJvLF72dhkrUy4XNpwr
KZp0mAogY9oB8sZebS1rsrAHPdlt9h/2RRGlUqfmiss5yp52wGoqZjIa3Z6Af/Jm
5TVGYh51OPRvSqyQ+3qtkf9VoAEBBJ4IJxVCvuqQS1FXhq2x1jRWRF7717X3MxaQ
+dRiw57jEXgxIOpq3gzbfNLmSdBpuJVavOVGN7gh4RTIkOGb1hhPTV1+6bC1U6Dn
uurLXN3pXuCyiHeXwrno/DcqZJjmI6vm+kNEMmHJSvo+ATWuGN+AiGHSQ5jQGILT
Tfu8Y4sbr+psyhgJvQdhImzJXz8dIJsrya+TpklYiCMY0ygSfKt1qabUlcUq6Ifh
A4s2pWjuDM39xG7N/nX/BMz6dMX/EUZypLeJFPn9ksMwYYdrNv24/lelA2XvWQVk
do+1FLZhsrI5PsuicdWD/wKKU69M8kSZoGstE5h8CpoVhjydu1ucOfNnbMOipu0I
nHf87NzBiTcAfVwWQKP3b94gTZbZwQj2k0z2PyBu6gyqhojlF7ntOuK+upGoQyE4
+2uQ3Ip1kMZg0JkkKzxHVVBt9MEi8Dn8qJXdIMr3HG+OGhTOp7UHCHw+bIPo01tG
mhfIu8U4SZp5TNimDi23VeNxDvQ+ef6TMnFKPUyHd2539jq0O54391GuPHjY6tVI
KOogF+QYdIsRjZXbygyDKpM0h3Pt+hdxzVOwTHzUnHs0wSU9ZhArLkBeLU+u5RiC
+qSFk5GSFAADLwu6rJC4kzKx4CH8HTa+N/2l9q8ov/cOZFbx5o3NnKPSsdCiSCXV
nXb/FimlZgzcxyo6AmJkPmxuRELkst+K1dfkiOluk8F+25DoYD17fS0KbpKUamOs
e8KkMraNIJZCO7WSLEWwL0kyyeAc8HfhZOANc4RQus8U7uhF1yE2xkGw49zY9uUG
r1O9rMxuGeIsxyb7M+l6GU2idhkMDrOPKCzhUn+USOM5dsumj191z5b3s55rL1Bk
XZu4L+M/In9RyJpJ7lib++KN3qW+O0b9xZRJOa815pRb2p2VWouWFYn48/dvI3Wa
moYnihBdPTEuwSt6rGSDUEaHIPJtriar5vh14C/6dbzAwYCZAPr3olBK/QEFrk50
4UU25kv1Ue0EVc+aBe7jSCDHF94iCPSXyORGP/YZ7eV+QAtXbOLgi4xxhwYco7Yz
8K2KnAAcdUQnTvEVe1kUmDlrTEesGkpUswAfmTMjEPnY9HK0upwz1IA3/u2xiRrH
xtZdQ5sYn6LtcuKR5qGNK2eFw6Sua6idvgqrr6pjxIK5gt20NO7DGFLy4OciGhxU
8ZZxqD4/+i19AtVvh5+lGzDksmfwHv2PkRIZ6mzDDDVGKlm0omIft6qZUMKGUlfe
b+ahDOb0WL/Gs8KxPGzVEQskuebrh2xV5ms5UD9XVj1g6i9rWS+pv+XAxLFXOd5/
+lNIbAZBfxnAYr9e1bcJ6rVDpKrxwE6bG/b6hgYMwu2/7Vggjvf6ZaLizxsJSrgR
BJ0vbG9zQjVDx+B+Hk6SvaiBDIpz/nJ7iJxRDJIwI5nq/5EKHzYm3AeMRGQgksrS
gMJrjhoQFCAU/Z5nOxnD0AVnvru9s46SbbPcCsNjjs5LToF8qaoG40nSbvPFRoDx
Q6TpqIXUZw37C77eGNp+GnKBX5N9CivfnFWR0GLtJCRdD+qBgfW4Ffg7wk0fqes4
PqlOCscK4Cou9IIvuHlKKre4JKy8WiFlzAWQ2FEB0HGSxXfad3zVtO8+JFFya5oV
g3kaJz4nXE5PqfWS5qhf/ZwD5RwnqM8Palx8r0MLwvr82K9uy7h4BAZGuCLm/zV2
4iAOXcHQRaookTZKRd2QO7E/t0n+UUuh2uWak0sZNx0vPMNUysmSFic51WNd4I0R
hKNXllBydAAhtbGyoFc8FLQQKmY+nwq6aXnlk12ofOgiZDX6I1MelMLEhEXB4GTp
uKHk0DjfAX4t7eo+e/ExzIJ2cc2OwlWghXz6vFTm1wIx8it84PNaXcTUJiHWl5zA
1uc5t97VRtRj0bsVNeqTUeIx/uzfCBV0kYCX/9uS10HAle47tieP9lzdXNIwtTC/
7QbBk2KflWX5k/96rdTieXIvF4aPr0OlWq9cTOQJqvrv0kiViiJ1wNZvP4FnagHl
gd2HomzbaI1Eb4wD1XfUOG3jZU2MJUuITxk+GZhy0DuqBPG+7zsknk0QZdpFSsQM
5Lj3aKMBEFyv8BFRh7Cp4WKERSJHD689v8F5KL8bm1JB+Xm9LrX0MhJdqX/O1Wfc
pclHYqnYLXqxbU11a2Winqnm36TJmY0+JWkJcR6JvFeX4eyr83AV63qj+cyO350R
9OGiex8zJJHP3JYXtJo1Y+TnmbwtX3mOIxOVCI5B/PSYUNfDqrRMvk8/2GoObtOl
SIFulfNkmz1OTkKdXZC7R+QgdfQKww2yyPKZTLzAfxM2LeWOaNZm62ZKUj49ocol
doxU3AUaJT6KFG4jxiq4aeLJvsDMA1/WUCrgD5vmTW7rn4gnhJed63m7pBxRxueL
6SaDKnmDMx1XkOC3HqetofXO7W7yu2mm29F4RK/d88mSOxlmtp46MZY9ygWg6RcM
CTFa2S0Gnao39oNn0i8ufqG/Thd7CSmXpzckWRO5KxMz9pMLKPqLGFV5KruTqTQY
LFZljOA0XE5TATAsxeVtl7v5q8l24M4+GW3dGswRj38iuSK6GpEQMszCxMJUKkLC
WhZ9013mqMGQ12LCbsnSrYG5vwrYbKRBbCLRt70egTGtNr2BK0QoDp5AWXvmLfAV
paZqSN11kapFtTYWHZ2kEC3U9IEcjeOGi8we8NRAQ0pcngyI5hNfBBtu5wExW0Q2
DvIyyGRL3AzrowsifaBAvpEBRloWY14LDtWeyc/zs44djb7Mbbg2LEdhYvUnSnWN
vieE2Z1eHJCYHldXks7z642KVe0CauuWu9T08gqkN7L31DoAh66fFfZGv8IX0em6
LXyg+WL5sBEzo2cC8SseqNa53LCAZpAgowM1mecxqJTGrOfMq0galkPxcZ45qgMH
eyqCD37zH/+OEolcLkM39Ov3zyXsLD5vpwOuZvP4Rgl1KDzFHseZxWjwg1tX3/+F
k5ieCLRj2ZStX/zWp6bdhW0uApqeWfF6KR8eY0rLK8rI7z18drSvnVaFXu/u2H7P
LCnrnCH7Ra+mMgWEbTQYD+del1m2E+PdtkpNYICIj3+YyAbR0c9jTeIImmnz49Cb
0t3/0//6crnH8P4T6eFxx3CD4wz8TK5JuqIPTUK/UvnMNyjebqdPKEkjIIz7JtMR
fNcELF9q9GbCx1YIX2xWBcmGFrwMbjweFljQ20eN00K0xcrWn50bPzhkujuY4prp
xnFLl5I5Z4zQGwKcjRbGplv967WJyUi7AC03DPBYZ8CBYv7v1zqdk1P+GzVEN84y
0mvyf4iWGZweqRjfl5WVu+J90pcNVXsnoAwkM0esn321JUiRUJSH58bts42hO+yT
ZHuWsIyeCNTDjWv2NozPLIWyybaY04lpfySOuWSglsitZB2C3WMmscs2uLlWmj1c
YsW3iQLNqzNyudR/hi+7zoiJhROMBjedcAjWIj4L1Q0udE0CDHLwerF8/iqNvJKc
oAyvCFKykNw9vhvWppaVVqevdI14rg60eElKMq3WvQ7wlUONJdbf1tu42VYOgith
hIBwGAPqhttSQqzj7VhXGlRoTYcHF0956RX1Y76OyTt6lJXHltf5CF4lixO07EiU
nIDDeEGaJpReBw/PcBvIKVGGwHe4rxEMH8KIT1amGZ9+AAh3JHTSE9Ko8GuBxNts
xAqoUHs/xLkh/GiV7kgLAcgtIVU7KyGav20uLGBZD2BKyyMqgbqzZW3CwU7MvnGb
ohB5OvDCrKMcl1vqkNnnnMod5qvBJvMmQSWzZKYpdxVxbWmBVhB7bAiCLJhWSK5t
gpOhBiCxgffNAMIlNU7GTzCQSX7TXi1tEwENoXVFSNRstoNibFchJgroy8Zr7c+f
TyuCD2l+P0Tse5tajdTjsV+t8wLjti1qrAtU6qP4QNSTlqQurgNsFduzLWKVJLkF
xF+KdbNJJN31enZw3fc2BzvE3yF5hJ+yIoWdOocyi+ZtPz83dkW693vQXFXiaaxf
S+Nmm30e3LAP7G6s93IaeVv+pthHhW+Oe7nMi1kdQ/MD2+2lPM0UFMTdti65qUtG
KdW0LBozVJUSOtP1tbarWCMomp1l7/ppBLghLO0Qgh8y1Csi65JYSfeqn37XeOrh
N6eWOw0eQDKpClqAxuXcFqzwLMoFDSZD5QHJ+Fj1DZT4yfb10VJZ21/tAJzu9Uwg
ikVJcoHLw3l2p1D2w04FKNx1IhPEyuJDGgR0xXvjZFbriY2YDJ4ZueJUzPHofFlj
sReEYntOAgQjgGPdGxi/e44o0wY+XlZ0/iJYKco7RsXWevdZ4F5GDTU0v8ojQQw3
JP+qsJ/Qzt4LfGcquMk0567t9H54AyCdIzHyCSt3mgr1Gxef02wjZvB/M8rBFULl
uVWgndnH724x9F5H/CAgcvFx6kQ1AYGzsjiIPxVZEJ7yWBiP2P1ziV9hj4vOMQ8v
FNDqkGNJf0S+5QaIY8PXB03QfX8euzaRIENzEAyNf9JRmNffQAs947nmFxTv9fRA
47SMR7GNtsbOKbRxkAUf9cHSe2A/qtid9c59OTvOnDoO4lodaVn+mpfqSWAXEG5Z
Z2/Kjl+S+Osx83y4mMBC9wdZC0yov5NRFsV5DFQv1VbDng/GijLky2UDdQBoDoZq
6xjy9neSQc7xonAT38RTgPY/Y0Z0LB9uR0gHzkkPBr9lkZaEOavLpo9m9FZGmevv
yMOnmTPgoFTt9r+1kiaHmTAGsz5JK97nFZekQDgH8PLWmL+O+2CbVrlzcr33Kn4e
9XCGsVDD3G/FHluOGqHPoJ4jmaC4obW33b4OKPgZf62S0dHuO0chyyH2nlP6NfsE
HZZC8OnQZOAry9GsS1UFgSY3ep2OHsojVyXbf6dHInv3vILwM2p42yehCMlhKoFi
kfLEF6hpcp04jZh75Gq2zguNKpgMOMUrwDs+7SsAV+mqusnW1KhG2zZd8F0NT/kU
1f1f5OEgEJeR5oPbtiumCTEFXcnY2DhcmHMXayrTp5IVWnRWBgw5czOtOE+jAIOY
yjvxHs3IAVP3LKzG3wiwGfTimVHZeWHdUSmZIyJBavOjrIZA6RMF0CTM8MT0wS5q
WOxHnM0UhDB/eAk6sMVlZszxJAlFATETMQakMnAVStEHUiPdwes9Vsi2shU0QRJc
LUWF/Zhkq30Ggsca0u4DsgZSsQ532hTEqowIkyylm8DRqVASJTJxeEy/fmdk+cvd
VwplcNDi0IDZ8yvqwWwZ3Ebgf+tXWYRSgZ1/wOuFfLQZoMmGV6Wegue8Zu6LuH8m
Ovl7UFCsfbbaROPGvGVuHuJ49aYUFl345jwNZpKRN17zPG5nWrKnFKCc+DEenMcW
CwC7QpApbF88mH7ZGC8tFfdY8bUGG3MS0LwuwVXdN7ORAd1y3sjKfyZ2ZChXj4fB
DXwVRGt2ybLjoTxcnGKftuQse5oChgPza77h/r3OUWe7rn96ydp6V4ltGCSr19dR
qaSz/n6xxo251Krc8RtVO9mqTUzrZlCHXxIZd/gSq4ri5gEB1CgL0UttLaRFzx/w
P/bWLyHMBDWeR4X0Uu7sose+kQqSOB7KLdZwL7y5PyduL4U8vw/GsAcrVSVVcJQe
jGIvOHm0KqjIzeAX3aXl9jm0bLmxfnzzRb8haR3BWd3QgBJ0+rhAM6VxNccfW/Qs
3mMS0XbqHkgRpIRDQ+ce+1a4mN/2nOy5X5wmsCfKF5WSfPGpMYYBTuJn/PoBmi/i
yoIL6/vxlin2j8sbzwK4eRbQsfCOw+SrKgMjvlSTsIlHz2mAy+hcsVcVtBb2gohx
ipYABzn9cI4OSZwOsgHMBb89ncTVV/QCio1RowiAE0jIF6jlmT/5kCcAssmXqnip
YmylcrEv54qzo6rwsvk19DV2lbMyic3BYrXcNQ48luftK3zwzTC55A0RDO94YTH0
/H5wl8pvEScd+wueRRJ6DUj6Ufvi1B8hcNDJbiMTHpESmL5aNENNB9aifJvJ6+eQ
SuqXsafeJEHCdHXPHu4UfkwGQTBaR6e5IOSptCrWOWK0UPWi2YDdSdAKWg8tD/W6
BNS2mssD2E0gI43YNBJoX0+CPJKv5RzpVwPTwHsvOZ8trEqh5zKRkihuErs2d0GJ
nR36A3oMdKwr+aO+hFhJQiSAIzYHz+AaJfYV6L2Yn3HvusJgrSjWCYJSKQnDCwgW
lqIDNTisvHhFxTQi7y4YcKUrTC4A+VsoEFd8EEXPIu9SmyBBKTMVDcbkLqMoVSvL
hJXP0xp1rpModlDITy+qrb1NQEb4UPEqnjxlhBox3uj179hU5HoSJPCrrJiPh7B7
sPZWJ1XOaB/96coz3/aFI8otpea0nDKdsEX34Kfi/FAcF12d/btqOxu1KxpHZ55/
aiorZy77po/XbJFRRADr/GQx0uaxHSinra2Al0XRnCI8/14xW8K85IPw0qQnP7R4
H+XIyo3YOWdWJuNvFvIl4SMgY4zfaYXr7KJbHE1ZbN5Js6F3Ob/0bddDW4r1pB8P
kcyHjn9q6fMgl/9trgL2i0+MYflEj1BHPYbtspK4F5aT3mXsVMPQpXAof5cmUmRy
wvoHUUAncx27CgYRYNr1Ev75kj8uHfKuFF9IZrj8QBIkEiFPevVqGoqRCXWQyJ/v
4YCsyFuMn2pCVO/OKKz5BU+w5rkEZBsU2rV9ldUsR4YQwRJ9gwBvstLggZHiwH3g
ceozz8TOLOSt3Dzrs62YUCIyoequ5rl+JDctCs4EFFtaNuYGWQ4/uKLaD6NgPHCz
xJm6i2HOukuJTgoR6bOe72k9Vu65Hi7Re2oWXwyg9+63KUXDVwtT9e+y6QiT1AXZ
keIIjm9VQWqCCZi9IH8IopOkt1PBNNMPY7YeGr2QoUGVgjW3SP5EF7nrpjz7ZmBt
3DGe/Hzn5eeFBWjMN4lLaIPjrDMQ8Iwhkqk8oZvBR1F6ZSHS5rykvRoetBSJR4uZ
om+I4ytzkvX22crEJun89iR08rUjx6QcZCdLW2dm/Nd0eghLWgkjbp4UGIugeJXk
Sp1B2ep7Ta25wpWMlMYOygTiklGktCxBUcvKVMzYH4eeZA50bZ8ZZvofdh4hUlIl
ZWol4NeOy6m/6soephfDCTW6I1GUEQNilpZd+x/VZyOGMruPCEGyYNpaizSo20Ya
T/OUIWIes+6a/DnYZ713Wm6H9bRHXjWBSG+jqRxeX3ShTgP+MLISCt65Ro0odxp8
92KVlhKO2Eg5vu93bHNvrpoIkXiyz3+HLwyBwS3Cll0DvJVAcVjCEo9y37J5Vxil
KNeGi4wDZ7n26DXnOzuEXE32r3oVYDPu5YS6cMeoJFe5XZ325PiMhlo6piA7yqhk
rTTaEjgGY9Ar7Yw31eIwdPaF5V4NKb3JfBWNZ/YsqlwoLiXog3Vaxgch2I12TZH7
kPnQf/e8z5b4OokFOyMZB9qU5yL8I4np2KpNREOWbaZw29j3PFxtr9/QcjeeEyHg
QgjommLp0S908BXkmsh1Px8jlMs/60bwAExp70iDs2FqmYNn0x+/v8SuQOjaXD9R
NDNSppeamU4oyC86dJJzIZGFygqKN38ril+ztVRwsdNk2886edhlgvSd6E2jIazN
jV+qsdzTgjfWgsKPX3o2EeYQ9rdePzqmxzDr0VIp1c9SnVI5tBvHu5qFTomWboEp
BQY+HSiSnNIY9zV9MjVszMJ63xtTgcEF55nBjDTtKA11HJfZsEh7efdCCpI6kCvC
XGsrWwwSssw7ptU93dqhCN7+OoLU3Dqcsir0r3BaoBTh4H5gdd9o7D2T9AMuRVRh
XCM7Q3rpF+HSh+qicH8jglH2DvM0Jz9ODbsDLb3StwPHmpjI22T093JeqG0ULG7M
dDVqM9+8hVVBkQHlBbHPP3QTGxRQGY5lQCowRGCEgTduLAFuEfLotpdnSBxnv8l+
ySZf2UyS7JL3TyyvLEhQJyoOwLRwQTa12ZcIAsmorzkG3/T4KPov7kBkoAXMaBsN
cmc91pChP6TfMlYW9F4xeKTfNA48ltQfXZ3SH8Hb79MX0B4zXB3IJqTDTioUA4yW
HQ3ip/UHpZq6iECdEM6fuQE7k+6cuZFcp3RmcJQYpAHKe65cXo5d7rLQ8RfibF+H
Xa+2fm2/NawOtnvhGQelr4w5vJgjK2IiwtreIHp2gIpvtyLA4cPw5V/Z12IUvmdo
ntm/yFQNFHILGL/1+74ti8sS9ENKgG1kDVZfUl2G4sbE4AkOYB8Q0u7yumCSDHab
hCZ8S44R4SSwlycAMxp7TtgXLLv3rnIdvRFFUdAgterRxIyBxdvC3JneUbsSwECI
GnGR4++WKiasIZw/JbyS7j3yTSZZO4FvedQBZ9II/WjsLSrkU7mJCFhPktz2gC9l
xoFKL80SEe19Qg/fdcRChKcM8iF4UJglae29gaKAULjV7Ok+Ox1ZHOpn2JAFH+cX
It/IleVIX5m0SYbsQC+rBDTQvFl3k6kkONY6itSI+mng7Al2rwreSaQjkUaV1gmv
28rjlHDvN7MCRR6qHFNCz4HakEOoqtIA05ccqkFQEftRmLqTkP1iQt+KOC4aFfu6
2aTr/Z2sEfeQRvzVz1r5tNJnBdJp8fIXnlrol3SxurwMOZfqkV1It0MmCvuRAY5K
liEZJAAYEceFKxkvR82qpg3QY3YpCHfVahKtKxM7tYTA3pTxhaXUOJslc9UXQyfC
pTuL3KxukGOnfVgDMXvekpwhvnpnUKbhloFNdRFGptFCXRzaUC1beTYC6wtU4L+B
OengfPW6GjEv7CM6uJgULSg0SvcMgCIEDZQbifT6iPjXouXdrKI8pTBfILjDOVaa
eBjPLn7JzSXvPWKwBL9GLoV9Ur8r6sr09ajVMJZJZNav6Llrr81LCJ3UbUwMYJc6
yGzfIcn7SHiP7JpyO6OAcOcvQg9XqrjwWYcNhLmY0jfSSopX+rf3Cv7nv0+HgZqY
xnJ52dQb5NWtolKVG1ebb24WNF1lYAL1XZarO7ROYwDwD0Awzx1f5MEfK7COZq8G
kh01LxwML1pw6C7Ly72R2NQpEXJUIhnaw7HIwneXIbGsqedpMv9FO4r3bOyRNhPr
lHrYSU9WIqtJqdMNB/oXwNwhDAO0jSaZa2eD/W2TJNS9YVLz5o9XXvAQOH+HKg6i
vFsQa/hFlb7ekiS8/v6k48e1YWqtgKEtB9kr6QLOo5RrwNov/C4QDblzAAqALsq1
TpEvPSUJOON/hSs9bzaIGUKngn9RaGDxvkqshZrjsRfjViZE75aDOeDnA0UAfRTB
8qq4qce+n85nZHXRm/BXiJp+jI8sFNrUY5/t15pTR2+uAzGC3mfP3rNazaelsCMd
WJ1Gj01XC9pOlwRm6FT28Z1Vea7NUkaAYH7GvC4XhbVzxWSR10BrnzTMHC5C4pdY
aollakaDQ7COuBTrEXQ6e4ASNFginw/BJatzH4l4qyW2sWYKjn5sxI7sG7TaU6q1
OmmwSKErUC/o3sLSuvSc5XpkoE+D6JsI3TaheDsZ4gcmaFOuVBSmHtL0H4lC8DHd
Z8sGH69FL3O25v45hUAQvbPcgAp+KI6efO/cnDPIKBFirBSQ/H+o9aq+Hyq6pq6D
ddnfOC8lIEXGkDoWHNTZD3Qes/G5qEFzuFAWN/yurg+4wdkl7E2ZLbSzB8yeRLNl
ZJNBhwYDCDsgeA1I2Atxe0sX+4UrTb5OiqjMm+fu9ZAWeua8N06pKDgpakapaUDp
xpza+WsD+g7hFS4yN3keoeySVqgbpgZqvgY0O8zRMYk293dTU4o1dJRnMZXEoq8/
s0hlx6YbHEe0txnvgLqPGM7VqzaGGOJA3/0InJvf4HwCmGKqJXeNZKy0wbxeE/tb
LyOsOrFBORTBMZSpRS3iz9AMuz1Dr4lJgXudAwb0Pa45kgwZOtayRto+B/zTu7DA
SjZ/U/oSDA0VG6TGlcQnn7jLjwlX0wf1z3nRNfaXtmGuVaD8LrLP70pjcaPJkpNi
4Xr3aIdzINczbD7rDRcteHyNpDkMVlB2WoSY0Kq9/OtClG4c3HsJjzTkpLdMTAmI
8xu3iS2XaMiqu6yX/VIohXpyJCSSj4eFeb9R4FFmX0DRLm6+miAjMXMyWcx97OO0
eeaEW/RmweB9bCqUoXXTp3eIMCux6te43qYyaAvHDtsK4B1i20qul/5rtKJCCqGZ
0LUPpd9q/+bNzsxj3FD71ftJKnaQoN+LN3KQvNvTge7NXWo5YLy83Tj16LF3h7W0
F5bij0jAfr0M2kfS6nhIlS9Awe2X5jRj/6gc5J+KT6Iy+SyXYZ3VyU+XjvyZIama
YS32QEZz/NuHARuqc3m1ZsypITSgli9NPNU8a2oJs1ciE+PyfUUtYJXIk7RxDAB4
194GLZkZ0qaXZlL5Ql3rNw+yTRfQtXYxIrU3a5y5xo2Enc6S+G4YJoK3POhTm443
sbiEn34qCill2PkiKwK50/o9LEFAJkA8+VO3s0WKNBJsqKw3E2abjnd55poavxD+
IQ/2JAqPbcgHAbdxPwq84RwY4yYzk7A7B85thecG22v786QciG27JSy9Ixw8lxt1
aNhxtdbJ1+KYAxHLGJB977cssAB4YzH/aGXHq1WEBFhNIvs6BsizzDvunJgCpHVr
FLNgLvXnAWEO9HPWsl8DPMUbrv2CsY2t0HRyg1lCoYkWNGDfKVBSpwlG59XPiURP
H7Q6IwMTWAcevI8BMH/DIzC9HXByQNVjBqb12lBL4HGv40TlP8YnhPI8k0/SFxcI
mpMQY4xjQJ9J2sdCk+L2lzyHzU8oWP6JFAnwVB3wZnHx10O5y80eMZ7cq+qcamuj
z7q8PQztMIbcW3gfqeDdGLzwdr3fCdvPi/8yQ7e9AgKkyXrxS7B0E+xKCU0+H5KO
5JsfIz0xoG/shB2bkDIfHra+UuuTG8rVkgc+a8wRn6S2eG0IIED8+hjdX0uin2GF
tHD1+ajdBKWem9KJO82Md2+uehb84POvNnpZxS8wnS5G+Ytqc//Nd3Zh7hsoZS27
3Ub8UHqKo66p01G6o66YUfMIUF2eIiaalgXx1OYLU2xy8fUH+csDUqbtPEbSPj6Z
5Gr7sglR99pbllX1Db3jYEn4f5KLmEf1iQA11pDdNMnNQLtCbG9kKljUCC59/J8C
8JeeWlugnqLMOqWCEjQASWKXRMzQrtwlC7U5I7g5P1TfczZCqFsCx6gcI7lew6lL
pz2IyZcMHUdtqMLCALxlD/Wh4SZ9o2QBQoNBKGbFN7L8wrZ/x1vXAlS+h1V8FE4e
r/t4wI5g4g8mljgrudW2x4Q2k+dEUjsnNJsJeZ1051kb8bMTEmmnfvfethZwPlGs
xPVaB22OrVs1adR0+lIXzZ/eZ4IlJwcVbeLRy+j+Dk2yL46A4Su14GBatD1xd87y
terixxJaBDCw/qJDhcj76P+/GuwvVg4PY/Ojdi+Lnd/v+Ub5R7yF+bJJVNi6KApt
uNn210lIYCa3ux3qEXI/nvNqpuGN/Q+qKaw9LXCjqEE6KNbA5Ywybdx6prUPxYP4
C3KimdN+Uzt7wIMNqsAMEwE0R4nr2WgYMOa3Q1GhIzQ49nUyQ0lQLd5tTWJLWveE
jb86Kc7HUAFYXg5TGGczQkE/A2Du/j0xGT7EwKc2QX88ZT2K3tLPyJziYslRtXEM
VQzBf9MxKPvI0gEtk6bmFb49tNghNLVeDPUnFJsMaPyv8q3sHC8Zn6NGkSdzfzox
q4Eys7XGQRtwQKGNlhnWGk+CEH7MYCsOy//WpYcdUCo24ielcJLTOheWBWxq0NCj
zWk1yJ/CUB4auvrIUXUDvrDB2nkoyGNBTdiZiwGQ8fV1mkbZTljMNFkfKCWRrPI7
mJiUkgtcZwETF1q7K9vzdPe3hWV8Ps31i2JCzwFtmoYOtZ/XC8/rirLX8wPbrnxr
MFDcOrY4FEOBZpJY0NfL5pzYdkrAhjIr7DoR3MEVbUHackerRSWmtJfaudNZqNOf
Os2QcvMx3LVP8CqcqMI2sGmHVj29rS4SS1n0amLKKW0yoorzO13Ls3m+LiwxbOs6
1MvNSCNPXanjhUHkPuuEblTZhS2CHfYiVnwkZarlHg4EhqNZjpXuyeZf7CBxrwzr
6UrTXYcFvmVGauqKwBOlX0or8LNqMiVyTYUhDr85OFyPKnpVBjWcKstJCJVSeQT8
Q8ghZ4F4CvdpMIyyYTlQKzx1g/thIqkNIFKK79UpcbvzPgiODI8QiyqbZgXmVjaC
g4WYAORjPjXy+W22rpy18Ug5UbfUEMdJn4nFwy9J+Iw+k1zShMfbPp8Gp2tdtfmX
omyYy8KEFiKnvxl/lUnog5yALDXgEQ0tsT+mEOTHpBUAgpfCqsgrrRkrfRzOVLhP
Qzk5hRksQ6jY5hOdIAb3tt1nVHS0xnLyaq+ikqq2yxX5RvpzOCsDPno/uPTBndGk
0wB+gw3M0zq9PTJ/Sy8RVUvMrnljGx0n/hh66DE6xF4KT9EbShX+/y65sQ4oJB2/
BwfsAb3UPRwVqmi5kSlwcahL1qNlJNNE0usqzC+6BDgrQqy0FK3GNcxKZOnCr2A4
B4dda701q5PiY5ymvDG594PKODXPnyFvoS/CGhyMwEx4yH2y4G7QkGNoES8afuoA
rODZ0B9XQdo4a1o+HId7DkObf7Nticsov291VwaL0WNI0I96fBEhI0arQpwwc6te
BJehsUfa0hPkYoWgwHt7cdFRJMa02zaY1EGHvshrgjGvUeBud5mkGJiRPfboEWi0
i/ymQp2P4KbTLFFaTrJ5Fu+fsmuMrjwXNkzU/mldZxYJRynqnb4X2lSFN+W7nMLy
AHl0xCY9o2DZx0pq7y1KEcsBr9WlePhI+6KC9trHykd7PzvEq1YJG/5p+A4FKsUd
xJ9P/SdAy4o7esElK2kpB3mT6CwpOAGdkobItClwJGxRI1NV/dmYVPTaO1s2Xkhr
LB0h+KUJkIwJM3F+CkSprxJvKA1JY0I7020lzSGSXv9NNQkIUWw4twZf0WOBQa4r
Yyo4NNnRWg3wcZM1IR2LhNL90ODCRcRF63KYx4bbbFFLSYS4b94dG75ax3Q6QFhs
A7Zg7swdk1DQsCo9qMjIH/A2olMVgTxWkHkfTbWEhRet+FuajLel+a1LpXAuuAmz
ouSDNV7rG6OxxCHKgjvDCakVe3BjDFd05Bl882mxT/WhW3w6sMpVSRYPbmSu80pi
aR7ZSTiP/SE/mallHpif7dcOixLeFGcL14EQlkLPMOouFBy5cas/zi9Xqicwyy5v
EJbisI9N7jIubhP3VRPqVGSVAl8j4Qk6zgYoh+yItupc2Zvx9KjWJJANP8rdB5c/
Sumv/1wVbfUTosvgWLS8HQj+4v2itZm+sQrt2QRLNLU3TcySDx6NTNZZoXNefgfN
nww72mH9A/4nVZ6/9WAIF7N63E7t+r0aYMDbcPSOej3YW3PUOUblRRgYvyChJgfo
wOFmTTmV1D0j2X7ol9sDN9/IDoTUc+AsD0r5pq506m+XLi1qR4gMNidfCQNvZ11c
Wr4yhNwyr0B2J4Gl20CouGg7TYKRvp+UMDxBXuTkEmyeIgsrSEYjG/wZl3HKd1GB
MNh5rTo/soVGnUgMcG+cDgoA0wR87Fiv72W4Fgb4OJ9XmHDfu2zHG8QbAPunl1Xn
SQSHGc8Op9Xx3A5tOQNps4yak0TwpmW9+ZQeno7OvW9M2ZCyGIlN2FYSlhNALsnt
wIGMr2wQBlLsawfFdN4nfw6Nw6svkqyjO4MCPs4rYE0SR8WAsLE7y6QgiU3iDB66
+tcKKeCoLvOlL8QJgD9GYM1vvsCidqXunyX4qKxp4ZzQAVG1KbW+WhlhkbZ3J19t
akkzk8ZknFoqjVSJy6OhvISUFWayonmQCIOsaTTe+kFfH66/BEA1ZwEjfykE7Bsd
n0VXbQZqTpiMNjxvmLjPNBQawaGRK1N2dcfIkqAG9t0Iyhr9Lcm4IutsTQ9oq+Yh
9IR1/eOsgVx02FD7Vsgrnv7CVh7zNIsz7mmxICgGG2S6mgrKYggUu4NEvXtwGGr7
/19rSvSH0c1chS5fEdcuTteKjCMiST5QL0Q5WMq/iyFNWxE/x5qKu9GasDY1MYLf
2NbSrFYbUnlkkHKoYqSpNBaqtJX8anzTI1wCfwXxJchsemSLXaFXYpzD5jnh9M2X
CIs0uAXZUCSRkC+B2hygsUQMW0u5CUV2Zm8IxJcoF0U2ODfRwBOwJWYvnjIusi1N
ITYUwJnJO36AZ/Ki+UUak21+h8j2DoFePtB8FfzA0cvNxcd7SbiGsQVpT98fN5Pz
c+pRNAm0sxZ7fFhOP/K0um2qaxruCxofMVjeB9Tvd93ceAu8/E1qtr4jETwR13ia
3SyMpwXC3+DuAGWjJo4vOo5gVLptcpoX3KScByfvNfZsPdhzjdzarR08ycZrOpq8
/Vsidp2/bLQVD1R7Q9sw4Qdsw6X7FYGq/m+YR79wveNibFLn8zFpmfeoP8lWVj8d
fcVvPVBe8Yh0+E/PWmSRmy4GJwWuUDGMZiEmS8n2pBqX2hETN5F3GvTEwX5ZqI0F
h5w6un0VtRlVy/SmV8LZdIfAhcCJVKc2Aa5TsKwpFgVjaL7jD4z3irT3+nVvw3fd
4g09gAQMDIvoX3eWBlLwdOzYJi9DJMJnfE+03vfjVvV1IQiGVJkXdrbORi6oxMG+
yWEZHuF9EsEDQNQYsVFwR73G3S7zCbriggi+WdqR/ICTQaBDyLyOFziphpOPWFRH
VdLpZU9N42hR0NsQ9xh/8f/zAD/PevAVNv5GFUGSMPbgzs+tSobhtQ6xJ2m4kBwZ
c8YfoCcaSOm4RBNZRnQyRqJ/Wu5M/f9I95sVYneprm/VZkXF7rALI8ZfqsRVY7SM
FNPWVXR+thp+NQqgyq7n1KK/kA5MYAjHTS88UBf6QIHPldgyrCkDxPB+VvqIor+T
2LrIzv89Swa7JrvX0OvcKKCX3r6J0j0K9zSOBrW5dDQ4kv6uTT/B7L9Kir1PjBdb
pVPHOH1eK0376EoX3U7ue5IxHI0CqaX+UPRQdypVI7Oi27IlzdXDdgiAkF3i3bST
88IWMjWk7dmIKFBwi9RTz8gGGXW200mR5C3r5dhNEA1bLYOxI7Rn+zeJn9CVp1Cy
QAIq2j/SKbl64sWG0ZMyt9vRU9/977Hnz273lI3wYIsPKLzcbd+IPTeiyahh0AbO
lyDxtEKxa8QDq25DDRNh8LOP+z8PXvziFKyB6z/QySZRcNyrMBQW+XCyAk4klf9n
RAY2WzSKyUQZr49IQ2iI1jLdZrB05kYhG0suI2A3zrs/GeB8Zv+oraMtNCmelNpY
x0IYqoVQRCvqhBdTXN6Tj1xoX9XpUFnkKQF/+zjpkjSBnp4Hq/+UY0dWKeiUX4GM
SmEsf9hPBGYcG7LzKGrn5JTkPkOV3KNOICnI7vOGao93+Ia+9qXlbi8if7kthkb4
WELaUuSEeKCnwVUFdeFblO5nVqS5SOmm2qQH3p6tR0T9sq7x38EoZj/cDq1dUnJB
KUqzKkxu5h1+N6kbioCUmEy21+/0Cwvjxr3erEuiy39iiqh1lBAE/eFzqQfoidaq
GC4RWCHBK29PwqUKpYAJ0m7Fqn9hRqsFa7GWD/HcsmbkGK/3PIxsAiQjOP/zCdhY
e6YbPYEUEYt6AfjH46CzzXcTPYSeYXPPXf2hXZZatYBUvxE4A4zmi2rUgHCsLc5u
+/7lAMwNKFWUFTBlxpJl0FCO0OE/gickjRSls316tSRl5niOZAfaSD9rP8msBEJA
IOMvuA+uSFzTghAXrTG2xLbMAJjp5BhwWPjz1n7ZvlWYp6Qz0VWxe4vyof5f1krk
kNKBiA8xL0IYDLGBrXVF0fWCbro95TbEcnAyShYQlRoNLX+PE4CIdlulSolNpNGz
7QOaGBUzbAUDnb3rM7e56z7QA4htQXCROPNNRRhPNyTHBLK6FQBr7sNnSDISYns3
kofbKUskyiGqh5qvvvhNIyfqvM2w7Z5oElnKRzoiULdpWFsx/uqxhiEJ5ctEjoJh
Mjar47o7SBBofdXhG8QnLz9Ux7jmUlC2mkngodhNPgFC0c7NeCJunO9YahqsfIcB
u5ubmVZyqHdg17boVTbwwqsNRWhdlhtUHExPWLfnJVJAQ1cG+iPkGZT4z/5E3BF1
JLiz9Q2M7ZSkyxtlAZxAZ1Fyr2rhswtLdyolT234MdkUjpv8MOck9wCARrCACIOK
UYpQo3dDPxsqhWc4iQvi2XtLTPdjsPIJuUtYPB1j/FJpJF1i37OZn5OiL80nXpRM
v05R/dJivli76r1lKSnQPqhTpL7n+rj8UGuZ0tkWIbcKDs7vaiCwg63Rq3Sqk+dc
8HvAt7GIKsLgPD+E2hxe8CjO74C2JyiBYOCnW9uziDMHVKC5cFO2zX6TmoYAYmls
KNUf7XYHjgMFsoHpNjJy+ZB0mt1xp3ide0otdSG6IELKOVgcFxemMgWEcljaPWnl
Lf1KTibE4w3hrkVP+5lrvtT4VieShc0Xa6bINPBwVIJQUUNKhk0aeCQk3AMyGntC
O4VvThJ0rAF1gLrTX/mOv9z4qvAgiDVSWs21ZdtXHF4Tvm6FNomt10nas36OKrWS
krksWVsFani9uXvn+5dbXo3JSuwW327Qt4Ppm00MPydvuhH9nKnQ1JzsPmtrMWuY
H0ZbIC3TLhVWYYb9nMhoKL2IepIFzB3z12Ok2L6+d2GjUj9JKBJHBQWpW0CaAR2F
QLZywiLPWfqWpIBTl0TCOO1lfFNIiUGsbdSE0xjCFussUnMul9JjOWEqjrGbab3C
vOtTb1fLlRV/vCpgGA65A+BObK8v7UR421nU4GML8UuIqFSKcztYVLjUkHbNJZE5
QWJY2Nvi+p5RRgF5Uk45eHLYQAA0BGOkXqrfNAPVVDYkgWe0zy9TsYQKBgn+QWcq
2aKkPy23Z1iYS3wOp7BB1wsOz2xKRNxF+2++TIZ2ws0SZy01brEEmGTohG1WbdPP
XJFR9K8NplZQAZ4GCs6UcuOq/5gc+eMopPYmtkndRhvMlw/GU7Mo3KpFRkDi2zcX
cYbHu0+XkI6T1ay1iVB9OimcmrUL4jxd78GDSv6yxQuOVSmz+74JqpFbbTJOj+9+
WXuQHCV6qG6b9xxXcNPwDL0biEsBDYe+9wCuDYEVfQQOrvn6/8iFPJnCBaTf67nc
rpSrbhNzSziwg46J66OZdEn2MJDTyw5k+IDt1TyXhAPHzUgxqNiMuRQNx9OZMWmd
Rf2j1+X39oHeUhhfeSLBPlbg7Epop73DMsaKnXCbHE3v43+Q/C/e0ApfaY5CYhEU
xxRcmKe6/aazddjscHEkXixJibMlL2Q4ZnsCYPC4s2XXrnJuy4MGTWIA7DZbK/s0
J6l6k4c8U0Llh5Cu/bamdwGMMsVVX4yBA7YSuxEjFkmGTAraLsCg9/VbtbMKbVfT
C5x2NrYrdYBWXpJwGiMXjrN49xk5Eudb02G5jK7m9unRoBRrrqUHSMO+Vd8XylWo
GmQplTMa+L5HxhbVDS5oRv0OAfmaAAPWJ+YXAnR2/otl2RFOR4b2tTzxY8O7S5sN
C5HXlE3y7+ZewocOFMrylPoyWQXcLO0KX4iJOLFZcAO8EJKqwp6QjC8PXd2yVw9C
/FnIqKePGXRoi54M+xTXSe6q9HRlTH4P+qEp+ebp/Tt/+HAIqIjkwliKPHIEDiTA
+GLVeVaQeyHxf6aC9XijUEZVl9kLqCG0bbT82hIhEmrUSYVNhrlHjR1wNVYYXzv0
d3jmMiWaB1Wa+CJ5QGSjiuprMVsC4mhKdQxYDFuDwhP9RUh8jPu1YSv2DpPRfPpk
aJIUgwy4k866nLNoz0WSvGUWqSZ9+Yv/Oi8ZfL+lvpNiCrm3UmkvcFIA/Xxdl3FA
jWnrQ3nNdgoXJyBauGooBTY14v5cGhLqwPU7nhd8KXeE71kAgGHYgh1S3OVjUK35
+bMES9r9FpP4kMFY/trd5rGe0RfxPHqCPU4hWuyrKu8AImlohacwfEFNzfmRJA4e
wVrUHWkRkEzf/lvyi5VOQBAfczES+iFfF5nd1LiL+v8X03YgVaZN6bs6YIW1sQ6Z
dXb9qPv50AkSoUTs/FjJaHFHYAdWbAbAjoQQeqqpOzee7bl4nKZ9pIuaA+wo4Fg7
SjehdWkbF0wnjwRwnJGsF1aER2i33iLm/ziTpFD9aYtph6z/a6Xt6W1MYPcRHJ5m
eLDMRa3O/CVA2K30Rkzi5yiVQbiEb0XmqBQIoK0u1ZxDMuNV6CO253DpQJkizQ92
7x/dikq1UZ0M9VSHXinWOnx42w8mvF1/6jY/NNSBisSA0tTbaOgyXzaQxeSGbsg2
8J/FaF0nhV0xN3OwcheD41iPL3EwyKP0q8HOCDVblBbi7K/2iVwOVkWvSvqXlV2O
xNLtddLpNiBaB3U5yqd0h768PIL7koDnmn2j45N5JYHnNTIRnsTMYY2GaoyG7afc
2OyJD4dMkIY1pY7/Y9pdai2wFLPaCt1/JwZZ55Fpz7bxY9fRpPGgaQ553u5ol65Z
q4G2T9hh//04IACAa+UkhPpNM3tRyjbCaAqKAioD5+kqBbuZ6QYXipMsGG41PSCH
cpYyGqGiV1v4bXDfjVgwTthQ715U9RMKfX9OnsqYcMumoF6djoa2irb0BO36lJec
OdBTlVZkFc4a1dRzPQ+oUsd/4YkmbQH9T0K+hFOT1JvRy9QCPpkBEzsZTvCsaUo/
OCUPXRks91S+Hat4Nq4jW6SQ4kG5FE0bClIBtu3RUbooMvoEwHh1tq90A84e8KjF
9a+kda4N2Vs/P2UQx8u0YCxs1SzouzTRni5yh6R7+/4J9/yNcRUY893sUmyfGvR8
lcMCv3azbWTcB1dK2/XTGF7ZCBJlUqyen8Mq1/Y//dhPhLs5i3cd83HxxJY8/AuS
4RXSQRD20xl5erv9zFn6D5SWgUgPleKfuwjzcLFqI6JZkw0SrO4KYLYsV5RIGaOm
mnbem/n/pUXlFMqwRofeue3MAdSRxUrYOPMcqSx5tC3UG5wsAEqqD7NAE0Rf8RPg
6Y9sqZPdOPPin6+XRSQAJ6Uck6mAgXjgGL1TMKRsSooeWbj27/Te8H9b60pKKZzB
WHLHuUxy8QO35XkfKR37IWkUQGVTtg0HWZpE48QQ7Ex52umjcSUDbT/qkfUWN4px
jnB8z4wyynigGyEt/1MmpAisZqmRycseNFMSuhVUb+cuLArDpHC6fXmoWhv78Dus
jALQVw+UhJnUyHjcyKNe0lU/az1lJ0m56bGrjL7eqR8OzXyUu/sW+YJWrLyfuic9
615LuVbnZuPHQa3qiJSOQRb1+Lf7JxfnQ8tIr2gTOkwzg0kbJMx/Hq6GwzsdYu2H
gKShA0egKeS/N9JlKJrWffllaBtoHoMnkeA5GdjD4OUP3VeBsLzhErzCZWXh93yY
2yLADLlQHHdYM1ljebln6UKP0iajgmssT63CPAHuW6K2jpiz4iebKVoctS5/7GiC
d612S0h40WOda+R6SthKq7fNsTQ1AZcKjKib7LIoi2Btls4SV3u54iPYAAkBohpJ
oDWN3QrSP6FTz/4vRDRCSv+TRa7l0OR1ZYRHR0TjV4z46CzCBvU67CN/gO25FtVk
d2OQNsDF1JIrT9cBDGbcRaVjjYFmIgk1Ct/RswZsrJUG4UpYpUAcpC1XgDaAXb+P
IROOlH+s/+4V7j/nBaakw3r8ZStMWNFkjINl8pZIMTDlc/SniLUIi07juROWf7Pf
dX/KQNwe+b7EHtTRwMvQv6aGnsUOCHG9MxZLfr+ewauoCYTihmv7C+E8CZYjLtno
0AlwM+wAOpcIh6ds8sEvJk8fAr4ALzazJTYFE7qYZmdy1uSflGjGPCon9rBA2DLV
9qiJjDoijCISvf82WpPNBBqp9Ym2RO1pOtte1yfJQQepFt5aRdZgqpT7oHDj0RbZ
aPRBkVbOBSm5YEGbsJCA2Gisd5wnpxBH2gkQlCC2EyG1Bsa+ZzHSkyRy8adR5oqA
PTSmWdBwutRikdQ5uZJEeeeDdwoD/pbDCfC2UYrpw6Ixw7pjSYxJLLHz6hr7/uc4
IYP5IAkIbR7mF4oLa7bdPIrKxxUSNqdO5zNuBgwxPnamlqHCNR4npfIXBltcqUFN
Bhv0Koq0K0V5v+yJT43+F45bvhguAFXzTwHdJxoy2YPZmDkrilJnNTzz4T08z5tP
oKV8fpuobfeHA0kabd3evpbELiCsrZj8yju+amVofWJBl0Wc4JtMzHNEVAEGSGhy
hu5WJ7n+KgdGX7x03F9yJDLUyHHPxNnK7niJgZN7cBx+Vb/wH9aLOyQF+XGDx4B4
wf7EkJAhUvE45e8jBnX5dpi4J5BhqAdN5S9imdt2Adp7YRdPwby5K9ctwSC5QUZC
/4/nlZrTzsTTIazEKAc/LHIc8OuxvRPcuapYO4Wts1R911P1sUJWCq3TMpI+EeT3
bq85kb8f4dZdVUcETmwfA1HPwCa8rnalQEWzc6uluTMmSV7P3bSK389KpfeRuirV
R1FxC4h+yFY/kDPos4hUelUe3pEd7kIj3C6dFDQ12m5xehkMGkbSoMJt9SDddSA3
Atm1oiGAUvuNOnQHfGKUe/5R+Br0fV04VlTuK6tnHtBxH5nAnUB9surGhbgAV+B1
t+/6hXrxuncTqzDLHgSw5rzK8cqBmnssr7LZH805y+YP0J/J1+3MkgSdZlwr3fmS
/UqndRkudRA3/2F/v8/JUDKOp4fO0J/nwl3MNkidCivST3EJKnmha7zFRybh2pTs
o0wTCTPWChD3HLGuVSPRxdIaXj2et/Ca/NXfq8fGaW/ZM02HCyVbkR3fDlappDlL
IOhFyUgGZkY8m561Brp7fZy4kyHVYTBPlJuGnIMihS6HkBMBmsYNaKW5rBSNMfP2
ClxtGN/1lWwFrZmiWIBvb5Cb0X/deyfWpxAT9wuecfKzKCIobvQ5IzeXXWUwp54U
bAHw8iKJAi8s4PkUEkdsmvPu1WIuVTTududEBkx7scQtztnY4BWnJ4kS0wZMq/LH
QrJHXu7UkVjcfN9Uzxz1gPpTzDuuLxjtD60vaJg9gvPe6lQXeE9NfTNYJlscpZhk
eY4KPfKnsLonyPNp27kbRIX4ixrhYX1nxfrfo/5SbDc7ToXGHW43xthLRGodFXaI
35pt63mIPzDUR4vK3lbv1xwN/Ol/oq81u0ZXHqtRfkvpVNjj3C+spy/dQJ25UO71
2lUuHu7d5fxvkYOZXE7kgd/OedpGDioUbRRudVnesvB9gHrw2a0fyc3sjsnfKAtp
1oZpqQoqarO5vy+xv7LX5TBZ/CfQ1+KihIzYxirwMWzzffCZK9JIZZZspkXlsgHo
Rb1QPZvEYqF6bd16t6EynPzhX4t9S5XEllBI8Ryrg7thUBbsVLAdQF+XuMrxVOX7
H+5UMeQTd0NVj+kmx4HiLqxSp0h6bjN1HDfR18dSy8hECk3a7VwKzCyBH0ZZDnWQ
/o6ENlyvATwhyu6g5trP6mE8bgTQ0DbKfxWt6OD+ei+ajY2HWy6SoYwXb/f87h1u
+KlP0YclG6suHml+EIaIgOX/zD9DYulcVfnwUsZet7tNN0wyZGlqET6jedowaJKy
u6mXONIITVcEsjy3udkguNO9qj3WkjkdI97Ua3wyowj8OkxXdWBCw453GzSP0FKc
+Gg/NHmEUoofovKiSJ1Ou7B2Gsq+o7dgYJ3Q5QaBKRJlMZjDpeIcb0xpZ2eaNcCJ
zM07y/dagqPE3OPU47u8jTqJw/zKFESq+B3aOk/HnmCd9ESKc3sOs8j1CAQ4d6PV
sLRBIRWR2eI/2do2OKEfKC2RZPinisXtTU6WAQJ3nLUWOtpSogM7ZAq1nNfe64cc
3pDyjMveCqOm2jXOTaZhN50tDL89Zx4y0+wzzL3Qey35TFbb2/geaL0lqzeU7Ymx
OX5HvgutpxNb4yG1+f7a5QEDRLb+ev9NnjH3Cla2S1Ylgj/aVFZLNKKaP09vddEO
XjaUqg6MMLsXYHXjf6n8jZy3GI7DzjjDJohEj6JBZzKHourJou5vVp//xAw9k4y1
6kJZ97WNrCd6Jd2b1mhK6nr7lpDNHE7vIIdQtz9VflzMgUTyxHsB0DwQp0OWmijE
HSM9ZO65mlT7JwhKWLtNewhdxeokHIHpfVtxSWzsHtuInSRW3P3PmPehUO/DSGyo
VMqXXn5adAQgN0sckmfWD4GMNaXaQt3EGUiiXn3FG6Nk8ZmEe/4d+ytFmZS8TMn/
6CMhAMwiApBl8E6EIY7sjFMB4yNE6b/9tAly8OQgex5tNhUfZSBA4lbdjM3aXJSL
qDaW2AthTniIcoQI8Q8PBJrpRDHuhgpBM2hSFPrt9/enIjDTsSrg4h2fyG8cwdOZ
iwzk0OIopA1CqmHtH1NxK31GLAnVl/rsG4ep+VgPizcg6yvsBJcqjPCG/09Olx8g
z14MKNasTBbxTNkxYa9aSPlnjEDzgWPIuTxW4OWpSFOEp7gA7+IGlGQjIJ9NpdSd
Hp+XoIk+trTDBFeLv5MO9DxykZv2zkFYUs96UlGYMowvU45t2D7dwDBZ7vumiJo9
hHLBDhFWKYRbz41PWIwmt656JP+3tismsPQDtPsmWXjR5vc+ugmYCvvG8baOi1pV
aqbAwt6sD8LZ3COqaiXIGB6iqINdx5ltzPX45g3tOR2hotEnkzLJ0h6RhA5Q4sXE
tfuk1ahj481KTBYNAyZ3MLutrZxAsjlG3g0uaJPzvqPd0xgr4ra3N/JBsF1aN5wX
oo3XFYhlEVadkwcFKpKT3UTmbw/b/H1/w9FBB4rkDN0iBt8CRb0tS4wx0IGL9gtT
sWrYfhTdgquWNIoUWS9bbTXZ2+WfrCBm/D57zGGi1oxYfHesRjXzjepFDcuBrpdu
frIzBNpa8MLW5voTFK3mezDWSvSLU7qolPjnH/Xx1nl7blGOsx46r1eAH27BoIjj
TXAXSczas66uKhkj0AIrJnVIVw7U21Y+aGWeCxAwg72tgZs6URxWMM6lfIuUoNWu
qLatB0pNy4Go28/dt9i0MYt242oKAvMZHMh7H8r182zdk1ey8LyHcPkazchK5Q1I
enajGq5sDGaxGJKs7yzZjNdflCcvsCUKczDLuPK02lKJjaoNMHS6qSzq2MXFRtTn
fFR06aN/KwyyFs9qUfB5tJ0qDRZmuOTmXVvrx/leV52gj5cNsrgPL2kUbpan2vJG
8U3dtUlamsyPkn9jiyWpTM/9EYSW4NcmK4F9c3H4ayWPuNCCk8g8MmIe6swo3QX7
tQOfuoXP1oGWjaE/kmlA6hkKvhFCH5DtjkovHyes8NORrnD9lNbPj46nLZFXn+Zp
n61laiWqkAy9wIhR8elA2WRqAJ1d0mSES8wE35GLcC6nW1o+hoN5HjpdYhjJIqDf
duLPddmKnHx8EUxJBXZY6ovb/CDcVgoFBMXYOzr/sqHZCwenVGY56QWEOswI+itn
wnyXOyBXnClRhEKcRuneIiJ3+PxqHt2m8SeWAfPdL+hrr24c8+VPSwHRhil6uTJ9
9vjX9gjMRVK+ss3o2ABc0iazDpOm2X4mcvqIphvMN15fgzpJz53dxJxRUtL+L91w
orJRBCUv+RYDcSmLDSi+TzrqNt12821WAhrbTZYTEzvlpryLvjxSM8PieBc38YE/
oetwgNnSIE1SN5xUWyzXspM9qimpl/OoiJMLoMuO3/mMXObu4D9hBUq3Scq0wUwr
5UC4D13hT2n7Ek2ttueefkdMMwYa6XdEYoksCeWy6LasBS0aHpfN2nNhIlrzfYJU
r8+Mn5BOeNT1BWixOMVC5Udeo5GbmaXCaOi/OYP+H5afDmTpUbYM6s63kawBRRUp
DtRN7RsNCimLFxJeytX51ssHbhJHqd7/jhrENl34kaMx0De38adoxCk5Uq4MCuIa
Nujqf26tbo5EQ9lT2eqdmnGbrIOdax4JdsBhsZLRRF2BkZlP/oAx4/2MNxTuGtPj
ZtCkq8e90jxZr2I31aSL5aqUz1qUuqM/Rm/G2YuBTgcNht5cNfkLcabgQmhm1o5O
KzSbMI6jg7ACTYzDJj85JX1aXsqLi3KLtitP5Qz4Z/Y3DF2/rPIlQXuWFL3jnmEP
Talft6JStxmg/7q97n4IbFqqfqpNYwFXEjp7zZsBH7Vn0lb0KFcoYNid6HdgEntm
Ro3UZDvnZ6wqlbXXzwC4MEKBOi99QeN+F7KyYn1LhQy8whRf6JgHjJxZC5NESFfH
8DFW4GfZr6v9P9kWD4127ZCGcrytEz1x3LWwoff20ES9qFgArY24+48t4GHnH+d2
lCAKgk+iGOy0+YExqyIm8PU3cFAglO/o76RsBGRR8lmd9ccBt31QQlcw37I+z8BN
EFU486JF9tfb/F2CBuSKwbAN2clLqFaapvAejUgyZqZGoa5gyKILRQ3jZWauOKQw
neDi8DFc3VwKj3MUrb58+5iIG0KqlaU+vpXxsMbkSc1GtyVx7FnZQsghkvXOY2jE
9uNa7MKdevuk9Jpt7+xBL+/s7P0QLf0GhjsQV850vc/cWUMeeuXXGCBZ7TFflzEE
jFvfJ2MWtWYzSAx0BeqDVd9H2/GubBRh5+JeSOM4qjaYtNGO6MqYvfO1xkE/ly4B
YuXZRTz6UI5D2r1w5MlyiFD5OxgUbJmhV7/lZ34s4eS/BjMznfDNnLv7gh+GBAL3
nC2ZB8lmTO3bn3NrVwz/bnJLMeUYXo3wRYXPI3yBK3oFxTlfr8ISE0+gPNa0e8yn
ktDJazlmJiEsktsMV/kYWI5qWKwFldi34FrMrcuFST8SQQsnJvqwrrAim4Wl3InS
WnoTDKTyigRyqNHWBudjM/4NLvRURMEHe1v4Blsaqq+edl5MFLcZ9Kn7piRDvw6B
VuWBxBmYWrW55URrjXGRpNRbmK6NiK3L0XzhMu6lAZzI+rqRvEDk0TNg0x24/X6z
KsIEy7S1C812n1B4GTzCnBRIV3dhz/sszV2r+53iWVE9Pr8kNFseBkl8LKhWNy/G
0e5N+G39cSOH1kKgod5aZfWtTEz5fdR78HOqPoVngJ8t6kgZNfpF7idvJjfDW45T
da8ZQwPTMOx9dfTc86prjCyZo6AMxs/L9nWuWdyyc+tsKJl460rlXuFrkXWL/ysh
u+6oJBmtJ45bP+opDUkr0ydD6O76KNzTYwzj0xsugbSsT2pdjREwxrQSlY2qY8GQ
0BCZRA3Pqgn+V1+luSGp7t/cYzq+rW9r376I+aBplOX32L4jTtXpak/tOc5GA6XI
wp187vY3i3Fx4cCciY/8RMxG5WkDDKjDEVih27RMWBM8I896LHytuhPQGfMIIDs1
rGm2txUwtNwJUYu4FwWQkHVwAvBBv6LkTRtP35iLhSh3vWYuyjs+5uyLvHcG6phK
yRqCqxteK380KoReshoPdj7fXbVuADqF/MXX/jcskZKIX7DUkHNIFWqdIp/V0J99
ZVQTPlc/YlobvfUi6bzblfHAlPLUAoUUC0yxQuEImy+uXTYRJES3XP5G8RCRXI4/
EMi/vZLqKuYdONJCSl53kdrXLk9rPo7qT0t5UrwzXiRbcEzYrYpaJNnhE5vdDpU0
uMJO54v6oKgmxW5I/Y0QArfoxS8XhtX6d8LsI6Sr4Ly8qnAe0/DZ3cVYnZal9QbT
kMUR37aDKzWHcoB5vj3VXjSG5lz82GjN7C7Y8SYWY+g3tAtREFLF2QBPENi45DUz
ZTnm839TyzHvCk4MvZP6PG3G19L7URehSlwq0SM6b+ddWl+U2BUj+2O4ev5GjeSB
WJQu4XhFg/RDfxkUIlz63oIq5HYlNz9gbeCfE/jL99XNXjFS/EykxR+LxTLnqae7
cKIeCFXVx4cnMbyRPkCaRBLu+llDOuuzIbJ0MU/H7t/91W2j5t07Ph3LcCKvcSf5
hDgKpCxtUaIPmHUZskXQhR99fGpEt2h/J8Yj2gprBhXlOfe/ZoujnweZy/JHuEWc
JWKXL+n2Y28ftLKq1S64Mw2mRtQNQPfGqnVVZqVtLWaBkshdGjYcVyxA/XIv9Ojk
9zs0FpQpNROZRr9vLQxuZF8mr1g6SiAFVTRpJzlW8zsEhlwr2s1FHgecsRS6d+bU
Qou1Xhg50CpAPP0PBDOhAB9rlYi1FyRriXrIeut5QnS7RprxlRAedifaJPeQ2QEQ
A/dvzyCMQ4arY4QWJ9MxtM5FdChZk8LBe0uyAEk/Wli+UUCZCZAC6Yhcb4F4TOby
7ZZ1pINVY81tQLjvSxzi7uH/S7K0cJkLJ5MDEAgpZdFJHywXpyWBEMRZ3T8nBBJq
413h5GnG1iaU4bBULgQEMk2SgknzQXmDZnUdKD7pwbHl0X1vgH/X2l4QDbAlL5X4
DyNwr3BYD90k05r88vBdOsoVMFyjDn+XJJidzizLY7xih8AM1knPjNjkh5+M1YgE
cjUR8S9HGP/ioGwFyJeblGQbqbKIvZtYkySOPg1/layynyd/D2jtmL5HAnPU1/1I
FoBup5gKTEfUCT74i3b9z3cU0arGTlib9hFG4ntd7M5qWN9t6aOHiHsGVfOgz9ab
NV+YSZpXMW1Vi/nas9CSx7W0ssCfBf3i5d6QzOPnbq+BZ7gDC32lYHPKQaK17pgg
h0699M/A3OT6FEgs3NG1G4r7iacCr5f15Ue/CUdzqFnRw1RJtcyX6vzMBnHJhazZ
TyVACvzGItka8YqPDpFm4zRE0O8c2H+1S4YNbjJCLAh9tIMoHDP1uMhMiinTn8L+
PmJa5Dk+qV9AonuMx3tubuVVKLvBw9b7N2n24PGcbM+6zqrE2Ibr1iSo5kPdEJWP
+pKxYABl4FX7fivzFdLxAC6LLGXIX1bHBaI3spZI5k7Nn7TdaW68IC2yB6S5abcB
YYrndMuU+/a1tnFFrDsN8wqqHsUqqQWWvpI1qCBKPW4lfS8Nf1YvE9/etDAyiVbW
qnHOHjgTr5rTGcqto3rqTMm51K/Gj/a9jGSoxPDBUYaHdw+M5mnztADg2+gUsGFg
JWrdlCDhVOZMQO54fd1vXgrIJvayRGSXEpFP96RIjwoeZfjymU/SBs9jToe8pETc
MW/Q9XHNKMP5g4W6FbRXa3hRO0FUdvWDoi6ifD6bnqK7qzeXoXeRshMqMcPKF67J
dzqyHwz5VGAT9LJwflSiucyQEsEoNHFbvgM+Kvuc4cV/HBWcJlF7sOcG06VC02W8
xM4J8hbdBqaSXmHEon3TbFAZzFyX9ibQ/iJR1KJUVCkvYYpwKRLhl5fu5Enki4Hi
MlumIY9EWDZjAruC/xQCET6l5bwv4MVHMSrsFdpbT0Lnahudo1GZT8AMbANER/P5
NvX56Dry/L7MvEiG86cwfBWcLwa0P0rT9Chc5vs2dY51W94sOJqpzjXqPASKmjz8
yvUaUrdPMFnmPJk2tBuZesiWz8uBpBkJ9Q+RCjwbl6jya0rQ03sDKdNfdtp5EGVq
huWdegy1nl6FOAXShbvhqaB1HyV3sX+xADs1PHG6wCl+xgfluSKqx36FzmcQWSxc
+gQXnBu72wdiNuhfajIDo/MdER7FUTCNB87Detb+AcW056PED/BVs800lDzGPIso
m/dXXVvDfpujBSH6szK1TjCxDnp6Z2c4O3afyzc6GiGsyzZkyN8PITQFQve3Sx9Y
mBa3TVBluF1h/FNvM6ICIjktzaP0VSrmQYLbmDgEgYbVsAjfASEU9muSyvt3ouQY
OdHUqROoAcNksMRHqx94yQpF5jvfd4N4KoiaNspBxPWqluAk8fPlfum/AZwU62NA
osdailpw0qpxexwwiEVkXxI7/zTv0iN3Oq3n/5NDZWldn+KIzP2nhJlaS5eBkhDc
48aBI7Xy1oZCrek7KqQHFmfDK27Eh93It/hIWTiI/gYaLQUp+61Uj5iuSmgr80eC
ZZuiTkIOJVU9kjvvlhhgnLV8wEJrRK5NKfsnqzeFuVyPqNeWFbvLkKcVkjzt7yox
SxIoAc98Ram0MKqF7Uuv1C9X4UIebVlIdUlWwCMV2y7c99q6AkaDuEn++Promv25
w0bVWaL4jqngDWS1+atR8gPzI8f2coB5IRfH0PNqe7sijWYWMeMf21SIVqu7OV9O
OJzDWNWD9OQnZIIK/5GwJ6672y+YRj7sWKRF2pK+2fYcLPlBsi6TV46PK5WV2P/l
yAqbaZtFkTAQ2JE19+qraRLjXzGeoJhjNy6iSocq1byoghbbWPSAHC2X5SizmQvc
3k5MxzHmkIUrNUhjdPX0Gog/JhQ7zj8yc5jRS77hMwP0T4xdkA7P+yKF6p61fMHy
+8FOM7Nj0AEQhtgxg4u3RaHg/NvpKy/Hy6x8/5jrDkWK7TQqQDCcIrExm44VBU43
pK1etF4Up7f4AGOxu432N7w0ZHAY5XbCXNnbgpOubb2SUkF1ZWgV87o4oznnKDf4
6MFzLiD8GMLKoSSFXBv9N7Ne8gdrc0Kt+6oKGEeVDo38isNNAE7vc4hErKIFO/F5
UyRYbRLgcy5f0mR0BGxawsGJ71Agr9XGBW6AJ+9Pejpb2ZmpIH/61LEZQ4GGtU5Y
nHN55HY0yOhLqNMWNF59LNZidB+htAJ9XTncqTLZ55ZBKbJqCKXHtQyRH7OsECTo
euWqGEsgEFhmga3d3S9RExS2+f0cnEhZ7aeoQ1Wew1cqGPXe7D275XDb3qULIRWv
thj8A+LyQYPhmB3gq3MTj5JstQucm6yn6tdOCH6lXvU97I6y8Qxzha9gns5JdpuP
IHnvvQutte+US5WKrehX5uLX9RgNwTxZ0amzKsq7+LF3Bg2DRN+jtMdYgxiLdKei
M5SjQb7rhbnctG9cBZ84z/gmyo85uwwO9rPYkn6+PYKpDw1cSNlxQqXHXN+/N+Ab
KsS60Vw07PoNRGPSnNcKk3JInH4F0LGYxIkuDCuF+4rgW4SckjZ6JLHzIED4+fcJ
8qMKgUWKX9yKmgonlCQHYiBK1W22BQJXaUWoKIU2XjDZojcTue9u2yy1iszU2Hfl
ugA/F7sn+9gttQ9q877Xq+91ZLy/d+vIXwCBfwy4deeEXpHcCp6M71MY/orCfaqB
IYiDXEI01l/yqjrKAVsZZOemNeV5ADdkPii19wmzk2dSFZ0FeyZixR6hdoufOv67
IrTiboy3lZX6DaloCaUkvNKhyn4/GNpjqOfBfm+Z5pERTROweuCDllOygOJu70BG
DHHtA95o5qBYugSWIF0ByBbHdk+qVx6S9bFdSHZ3CdhnKoMaYnDoS9YwGMZHzrRY
KQPYRglfnCrbWWP1tp/s1aanl7KrS6tXcNI86+JwyM/EYuKhTJHtL+vqar6qHwNx
3igIeslKovmCd7V22b3J2ohJozZrIwXMpmDoimRGxKQl4E+erRWoeubMypiZ9LGR
gvwnHbeAArRMF6WfJLZLstXlsohDsjhqrv6XT07jiujM+OVO7xd7jTn6Ovtzutww
L0npl/cBz/NydhWeKLQUwsfchKl+FAgSvjROel7Kk0Hxk6guH3jlkQlh4L+Gt7ki
zIqRBQ9F4yj3JKehH2s66LIkjBNrb2q1N9gjcYY+JKgdDRr5uvCGw0D2tbyFVi/D
+WSzlVYMILxHbHcj+A+t/sJNORIHDy+2bdMqFTlS8N9BuUI4zaQthQH0mp5XJavD
YtnM8ePRm62CnOFmZlJopBI97acUmgy+vTzsIo+PBhv9U+mYSYiw6JPzfMyPow7O
iI1BdfBSSXuRkKsdfIrDNlL3bEcKcvWy9MUcVGGiLcm3rQ9hRSvFP88iXyfzCITA
DCjdf4IX5JqlwwY5ry5RCR56pfKXREnERY0sObP8PHWtLakrFhYzKQj5w9+0a0HO
KBmn92Za8jYfFkroLbA+gkmNvN2iTPyTz1qEJ32atASP+V+KJKqwtetCUX3MrpcB
3GkiHYnCQC67aL3ixxOrpOJ63Czx/tOhzHcRv93rPiUVxXUYHXMXgBvgspZ6ydBe
Zbg4il00dLidXvjRhhcUm/6Ju6neDNjQJ9oua7azxoPND0hjk377UnJw2JE4BHex
ND/OPE6XplxsG9Y0mJAJMg5iaC+5EQ/SNlXIeV0GcyvHXHkmAXzrFn7cEIY6jeBQ
5edMNkL5L+4lnvoXzHoB9pXNtcxwLo/TAVzEoCquA+6tYx0S37TWbhi0yJWJI35o
xblmbnev+vSXAIz4CJG+RpXtBIhIWeRFsy9hSAY9WVuiVjVayZelhum1U/ZW9Wj6
DOSoMWf9wblCPd20OhJnrxceFygT0NgC4YLRklCPz7BkuDBcqnGK32Okbw/0RaEL
49EAEFqwCN6cHFEMNVjkiS69hiEzlrUKt4cf7ygP31vwe6oSftiG52fgOB9ut7N/
pah/vk8a/zzyMU5TiA8bP/hrioSNthgFxht5fPKH4G9n/pLykHG18H096FfyWBBO
i1alAhHvKo+YLh/vK8jtaSCUiicizF87aDHLryvQHs+Y+MQFAHa6KdCf3/BS4YRs
Gd6lcfm0jUALI6aR99rCoSoaqJIbs/Iw3DIxEex8pCJiQQq+qxaqNH1u0Sek81iy
JFlsUoQO5AakE721S7oLmA3FhkL6zE4yZ/Fxt8NrZSuSH1804bgW/SgIPKslcW0a
BTM7R+SW8vcGPqn8ejWy1pSCygQQ6GCIUjQYR7ZwclHPx2ivQGYgDA82Tn8UkHov
Nm6mt+Ah4nX3LdZa/p7u/9IosJ4jcWFe+6iTHwi3bNGDwrnjrKo4xMEoXsH+DrFb
uK/bcPgipU687Co0SR5HMZZoTp7Pfs+uARdjy20ULWPXR95WJbv13ab5w12wG7LT
f9X7lA2bAhrfwoaPWe6KIgWIfXQuebMCyIDFVYff84OWfV1AiOl+NSRY1+RS/6Rq
zjn+Oip6+UxMm44HFXak9L1zvr6KpfYKgDvsOecVHdiOcvEoI2mZdikUft4x++Y6
2mcOVqPDjr7LRq1MKYJRn17w8sq4zk7G+3AbqiS29IkQCAMmmmGWJgqzw/lVT0SL
Gdi05G8iyAC6ntQFPpenG+cB//akiV6CVYPRlCoYJTIP+PRcTEVhVho42zJLGZ4B
x/qzV7LlXNidWfKBxhkZNEHdG9PIHamzzUDx6jr518TP1AcvheLKnVLH0wdMBWUU
Y65Ms3Paaaq4Xu8CPPk/6brl0FDP1l0ZKDMJo9Db+IN/pmBX3pIqryjKZHr70KAZ
kIj6Hfm66Mnx3rrskUFKQbmx7SscLWA8OUSfUVnLogvhT/Ikk4KBIy2xQRfZcnRG
y/tIPMDGiB3U8kK0isuNpyNkuMQ7ZXB/wcpxYw0haqx/5ZrIX+p8y5O25wKGzks9
ffQqBO+vo48g/w9xneUOvCjGixWrPJ/cnuhDDP7f7HdnPZ5X2z3+eQ2njocDj8fO
KMM3EYiIrdK/ye8Jaic3SYRVDsuo/HkNIxebLyyrOO/omTHd+TH+FOcVsG6+eT1U
QXDH04mImXcSaDsyIq3BlzvtDAIXyHxq7Tfz8NhTDiABLo0uLlCAdQpJAN0B5WpT
bzd3aFj0kG90v0iTXjnQqD8esIrFZ4RqHBHoifdGbItlO4Pd7QZm8hkPtiUKvPWq
uBZ5zBwnfJ6mWC6EVAbw6U+4bB/jLw53xXBfs4SXZnusZx58+XHgL+tH5GiGoSsb
GHU6oAWZSujGvgDuhs7xkazALkAOzFag5s6MzCQ+Lzoy4fKHv85vT1NYKXL/KpGx
XmbqQwqvmRwg31++UMNw1AmUBiKTif9Tz1XCQ5T9AIMnnKAyBf7mwM//6RBruN8R
FuzhjZ6OZJjD7E/dhpNDsPaFhOfWZ5Acy8INgNomKKTQ33Xuq3nH0McUpOQues8q
rloyD7QF/d0j0UAOtlIlebhwx1w+RXe6fVk8X8YhJDE42GK/bnvS/wtfJ9dj734D
WOypteOEcDQw97lv2C4iaVDSx6FIkt+2NiK0t/LSvUsbyo59ZlQV+zR1hrjbWxVd
vY+dAjz9mWiUtXW0z2fWdDyuwY13CPiDzhu71xbdPtnbpmt0NvEP4XeE78apqzju
HNDgfb2jJQJd2Wkrukyt4U8rukh03G8yAQrJEb8DI+EWsP/eogOecmaS6ejfEIca
ivmq3zAlc0dR6uyPkLokyEeRifzPXDproriB6s61GqrQ/iDvDTbAXBxRK/8V+LrU
ZkLX0ytYY4TzAPrwHYFucpReUKipja21wO9rxh2EYgxSOEqddSVDloxE/O4/eqj5
9PCw6mP7kcuBvr1aE1CxIZ9oWxtMPrQjx3H0Ad8HgjX/4z8TJyE3x1o5g+n5sAiv
QEuYOMd1KzIFodfB2/idxy1WwiBhSfHy7zi2eqDLmz/zusCr2Q50cfjsxQzehMOU
PBEEQKUJ5ztCww6XaT4L8kL4lAiHEo+r/qfhBPvZ7OC+/mP1+5VZCc9UxuD/eTIx
0Qj3piCAW/35DcqHh4nLZIVix1MzX26POByMYi1TkkgsJoi7EnSsianLeDELBy/z
EbS7vb1nOqmCvIGRO04WelpilaPsPpsrsz/75NrFCXjSYtLHQi3Wz04uTp3LtNRy
sbcYWfvrWxWu7JiWPN8QZs7cVKsSdulEEviH/1lJO8dx96k5QI0n1veM53y3FGIU
X+wsnc3VsjfWLZN2TRrySaHvTUn1cYTfx7LI7E600ye/cq51a3/906AB9Ew6RJY0
iZlp4HvN8Ajn1u5XFcWiDwpRxySxEyHd0Tvp7QYJtuJ493SDmanyaMSQ6gUtTsCJ
mdCY4WO/wxEfi/mkByTFq4GRbJcMYtX8iHQOf+3GSqzRFjYwRAh908xIn/I4WQYY
X3C9KtbCmQmwusmEqU9MEiwz/O7oj/3R9WgGXBjkHKikVli7+CjV0J72fYA3joQZ
G7kcpbFiN5crN1Uq+g0GjZVWyrWRgy1GE/z+8wrNFTR3f67vCE8zA4zTfofoZdOc
EldamWH3IsM6xobd2o9JtNeYossT3pNG49IQncsNy74=
//pragma protect end_data_block
//pragma protect digest_block
2HBuU/n4aRFt8Ytp8d5hR8qUSwc=
//pragma protect end_digest_block
//pragma protect end_protected
