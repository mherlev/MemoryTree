// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:47 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
DTFWbtFythbPuRyD99bTRnbItiUBt+F8wD0o+7RtbLw7Zjymq52RmcRC5pBFtPLw
5Xbhz5tC19PjGUVXtL+QXk9HSd/56e1a/PDQ1XFhYDt2H0Xd7kHxwqRys+VO5jBj
sLZrep5fi71O0jAnyWJPywzImWeXHQlgZxU+WBExCec=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12448)
XpQs0NR5ZXB6MUMoFtSZzS7Caf9zhqq32f5axN98BEqvTpgrEsyAde3DLblkpCmL
6FpMQPktvOxFnfzU+byclG8H2fMZ1dEkM5FErUinJN/JnsQTMEzf+8YMkOB8qvYd
heFwvxfD7FxYf9avEqn+RS3f+Jk9s/2xaLBBObbc67c24d7gYwbG9LUieTHmuZjB
q58J/NM91QQPYKJbRC31s+uIxBO8lBkLsBAlctPPeEMYImHq5dDGedxp9gg+aWD/
l1cV0mM2592HsQXBjjExZwGNWQRIyhTW9VSDZgRWPYDCkDYMiAX3WBeKRExv0Kny
nJKV5oT6hqPXku1Bh823pSjdqwL6PPXJEkkYFhJNOtZd1SWmJndhtO5FK+F6U7iC
9Fa3144967g33PGBT3PeaoOkZSu6EgMllZ2kLni4RSkFxlzJ9CwIPeANhMoY27HX
mc62y9hkwRwLkZD0NM1CRAoEVpOjDiMnjwqLI3ZJhD+Ra6JDM4c0DK/qvFYMr7HQ
B1xqCygPTdFlYZc51yxWqO9nwTGFrlBMZ9dcZUFIgn9OqXyhgpNH94AdV4Grs+Sm
w8fGE+BwO3lr25uhjaaAQFXaeu2CyOslILSK9FNbJRQ8mYKYA1AQqkJsEF7KShRI
oFNgeT5goUSY02AaFw+BQ157hnKFPedZ3weyvfap8iq0ndbFF0bFF6mKV8UyDoP0
jIDjomwqn0Q8cgFLYoB504g8yM6WLmZUK2JM7+Is1FbtAl4ldn6Hw7DMi2VJeZta
dbl3hqJ85CtJCixg2kF5zZNjol5rj+Tj5Bx8DTbFn7KXzM2Ozrt1NEHD+sADAjvI
YTl4eBo+DpHYrG4Y6JsB8/ZI9b3kaObE5Z7JM2WWH5btrcjJfo2QeN9Q9iIj9HLd
I9JZLNWfX/IS/B7oIn03sven2m4kfbeZ3J+f2XKYOn1H04haPgN/nRi8ymr6tMTl
aVOTj3bka3AkrEUXsgfX2F4ckaLmpj0waf2eaSZYZnSNqSG1u21isV6sKakqYUU0
tW5H85xmYCjtTWQv9KDSNfot8u74Rp1SOuJYLdXxD9kONTHr66/PkZNoR7jYTJJx
5leH79kVG4en2smz3Vycteq9pJ90dwD+Yi6DGNVZHKDQw2e2Xr/8uecsuaTHlrjC
HeAFwvt6exb3kTLGZDX4GKRoSP7SK5Ihk4ZsM2yFKE3SMJoZgr38fA5l4c6wVjQC
/F/D6mjhjgS0WjPqRzNELiSXgv7f8grk3nF0wBWuB4Qppp8tsLugncGqqguYro/0
aqfiiRhdBvajFRv/V/iPO80W1umO9Q61HokvIEeosza8yjcKOykrprNBfA74+Bj1
uU2n4ZB7F7yyeGurF2LvJ1mMmRbtV9qSY+28FOeq1nbEiVh3ddeIQyol7kgUajsk
iJYPU8qC2aqlCh9XDZQxUcDv4u3V9NeU5W9L/YUx50sZ5CYNJometzTc2MW6iVYe
+w9InpybmOG3FPoO9ZDpiEmgRrX5GGUIBQdmRSwRWQjfRpBsUjoMhD28VhmItYSl
TP7FrRB6V1pJ3mvGKXAMdMOQGHFBjTQ1VYBsdQ2u2kcbEmVtKvAVRUTOCGmWrs7s
lV/tEHiWW8AGs3hNl0Df1rN9/bB1juXrtd470LAaBRrcc/Ybs1JcFHIf+0lxlRA0
jtJrqxMDD0xYgQlD7Rjy+CVYod/5qEcZfX60uSmna+GiESN4AD+9fx6BWDu2o9SV
MNMt+wbKf/rvWfQMTn4/o5ZTW5uT5qOpbdZYnApG6ir3I8Dov4t6y2PUjsWA0fq7
uSm4R9zZ9gPopjOOI41JjZFNoubepfiPCT/mbbX7HwrejdmORc5kvLpJqvVFpASn
lnkYP3XVOq6/rQ9JdzTh/voRsvjdfBiZYdss4DX2g3mNhnbiW23rqFtgA8yM/KRB
+ZmjQLOahppkKqG4W04Tt4mXi0ZwR59BlBq7RZYeVeNvIRLnVksZhnqkQYq05zVO
c8eBkIJzmi4oJMU9hlpJ+TFdHv6Z5IfKKMLWQmrNNXNHIGVMIyCw6qvvqj8zyt5D
wd/eIbWbxpSvBdS7QkINxqeNFxTOvG8nTyWAp4m3PF4/G1Za3KtB5LBOFAkvT6Ym
yjhzEIn1v5tVK3WzuBt8qI/C5ADZRcoLIBMn888BMsGbi7XQgUvhQbU5oOeFBpM3
SWNPNeAhsLi7xq6L4ZhLKugwjPm7SQqIsCHjglDycuvG0HyGPqmU0oi8Dtqzf0il
tgVcoEelBzDHMKYuV7x2n7tg/SNUN7qbYhJ0wV+GyKRrRE/3CVYsKdLr+vD2H1H5
NB/yab81a0RT6kWqIx7+ZjH04Do7RMvXujZLj6aGB5t/gR1tRzdXUfm4gunzJ7zz
j8XiwOVJxF/q12YTYo8Iw9iIReHz3r0Sx+UaNN1vDot90VwvHip/VH9ATXazmZSt
M7pFx7DgeshHzCsYqqdfPcQlIwu9RsJQQCSpAHI03EesxF53OrZYdbVLtzhDWCPQ
+E8Ug4QdqvGolE49uUI9o6hYGWV7O/TIrY3kZ0v9tpGAekX8ZNadIjyR+non/116
S+CvkJn58RcYZDlAqGpDXnSjf7vKgh27uwOnZ12Kpwtsj98KWmOwwhO1wfonrcoC
q6S4N4G0w6HXGnMXwuq1B6k4uF9wH9kUfHBQ/8yntfPO/XvUa6GAhzChuj84Klls
1RcfDze4Z6A8Z1sH5/IPx6yf/00ZWE/8h5OlGjQM/3+2PtTgo13ClIwMDsfN+2gZ
k5z4d+jW5U7W0KnNv23SQWrnUMF3Mgz34HGizH89b/XzSytjsGFmz3cWxixka5zd
xDebpLbliDkfCLhtlpLeETImFbBesqfMKYOefuGhrvaYeFKBdI7VqK1EGJ6JeWKg
6rYsN4LrV0oGxIPbkQv5wrxrYX5sd3kbzNxtfgjRX/4tNk+0BRAnEO59jqRUYlcR
23YTR8JU3S3ezfZ93gOP/FKExYoV0iliIIXqfUz5H9hCGoG+FdYVKzTJis1b2vhx
Z+kM79ZRYS9RggaJk3NbEE8rt8ZnbtLpmWGbGcdlPSEF5d4/EcavgJ4b0/MtnI6e
lTjI+keOtKw36Uu1gRpoO5Jf7VGJoEDlq5AYfNwbPjAMFl266rQDaokvc+1PmI3A
jkFI+SnJdEzRxhcMRWaz269hWmPFdQZWK88xlo7ADhL1OmO3icANS+SyvMZte0Ah
EhmCfFHk9ptA6nCaZkdeVR7ebfJX6FcP93mjnbjK9HiNgywvNIittkxWzKpnW7Sy
13G/yRAvFmHV56u8cfNrZT+n4OjBVLGnzTdT+xmhW840n4C4q3INOU5hwuWxmWmB
ruSIvRcwGGYWlIZdjDowiGbaePQwu5ffuTzNmXCOTo3nLo+h+wBTggpGwG3V1rPQ
JI6DWe7JrkqaUlVWWzDHlDXZ+l7Xd2T8nR/1VnFfA9hVU3aNlecri6ZSTAqRxJ2V
epjbVHSgGgsm+Mt+2OgEj+dqckbVMYxwIg9M+fjydLOi2NeH4s9iUQBbquQPUC5X
bMd0hyvyfOy9aHOwrgZLMrr4Mw4sCFQR2PNJiLdPBbz/Egd+k9cTS3tgfoT64bC+
xnOG05gfTWQGoETLHKVq66JoHcb5bohRAsLbr3bVYCmoUBGD+SLU7IDczWsWijHD
ljRQO72GHXPyU6FCKh+hXmuLCan7RyQNZd5Oe+Di/4xzOdslTv7pUsBqfYFdhJBB
CGX/xPH/RdJXcCMbyuqxCp+q3Rg0wN7sDBQgAPlbKxPQ6aGuybeFXxqZaZS8tkih
hU8hZhfxIcYw1LKrNmLeHbB15xOo+2MzhE/Q+P+JtVX8NmrccrvidBQXsZezicCI
jKtrEdJyi/1nUYskUXSrgjXPU8cRt3qnNd9wlcJDiS0dbMdY28/Qna8p+zx3CqRk
dckYdZVJOGfizMJFow6VOoVeC33KC4EPuOqX/0Vue7e5mznEXIwuX0WHTMN5R+E2
kOSRuk7FMEgZJPxOldznhvok4fPh9Z4+i75IngTmyOaXzrpwvjh/I8VRF/gDRXra
EVfGvI7k65fIzpVt+SAkkMxtY+WqVtlwXLE8cHpUiF+AZeB18s5XB65HBPsFbunh
x80ob9TYj9aT1NZcD5Z6BPJsN+4h5tBxW6YbpvMIzTwzmDesW5Cg7QiOUshShRK4
Lc1FlCVJ2DIDWdKYxKvZQ7JTjbNGlZ+JArKSIHg0m7gSkVX6gOmI0lBa4ucfOQtF
L8ItOwBN6T8tFEcZ8cU3tIbaaVk7NqTtP0+T2O+wN5RNUYPc6AdUbocA/yON4P3N
HxGKxWHPFzbu9OjidxJVwDyft62Bt9qhe8k5zuWHSmuDFBtDLMskkBhia2w5BbK1
4Op8o3kzU9to/vPDtNC+QzbDYVy2f9CdOJ6vU/0OOyY9JbMKiiPHDa5cHTEfkFSw
C+9GJZG8tl7VUswULcOLxcd9a5E0PSlquGCHGIS0kMe076pToy/kBhmS5CAVid+u
UmNlXahbQiJ3ANXs0eHlaJAPbYSGulcYbHTfoqluJCDsh5rEjYBMkrlDNg1smduL
KaX+0vnRBQ9yD6Y0S4vLdIo6fSlsquDZr/5OjO//56Vds2PE0IORI2wkBmzhjHJk
oiFRwtSjFpH9D8KVoHOseGO7poIZFutrexFyjJL1jtcjGOWWOkbu6t3RKfuaOjcS
NBqAcxlAO8dCkR4BMWFxRC6VPBHuMrAHDuwwgQUJ1bAZh4dtX7bRYp+6J/aEg/27
T8KFKUvqynZ/XbcBH690xrHFp+WaL5u/nrvQXWmW1gFnFX8FmvkUnxgg7jf+jg+O
P7Anm/OVms7s6usVwhrdYBH+KQc7xsOf2cP2XLSXvtL2t14dejZFbkwofkiDs9md
JqNJW2Eq/jDrIJO79nxvrxjffF+n6MUdz6weOPOAst1Ht8Lr9uj/6Els3JfGWBUn
E7R1gcQEcYz9hACwQZwSDdLR5uPElcYFleWkkqUN1de5ZysjzCvgZEUopE8/37RB
iQo+1Doj8+3966MiU7nHK1XYci1tehYZM9juFI2qJvdK0c4xFWKfeaRuecg+Yxt3
sR3/nSkYjZFZrfeR1WG2+4JSkFo3jgrl1E1JCyg0j3xdq+to1oedQtbQuzDHOH2h
K0XikXNrDdzkQzKwGG0FK7mC7mO7zoREshT5jzD949Kx48MLZD9VQXtzXk0Uu+jG
d8YTwYqC9bnaV9Mk15zdYzmd2lX2LTjCbvr4C/YdMT37dtflsazPcpXNXG/FJVZD
TOVrqvQviMrHgKoTOc/I0SKECNpVdyU1LjrysFvQtCFiiu9OIVV94rt9e68YyQk4
Mw3r6bwMTqzqFMlKlOKzkhuORybFy57H9J8jELi7lOg+lIjcBsLVQjpy0kOiMg4H
ue7u7MblTdI2moEHcO1wNSyuVgZxe0o/lV60yA1EZUHwzs3auQKKcpg2tR+q6/t5
XM9hjAg6ezmYPt4bXmSorAqhDnLATYldm9pHB0RrKH1v8BFl1XJF5mzmtE0t2S+P
U/0A1N+jYLFaOAEUV/wO5qDOO7ZD0R4lXirklrtoq+oheC/prYrLQPT/ndo4YhiC
59nEm8nMg5y6UsZzCVoCG5q+qKdYR/LvyrKHxun4UL0mWKbU4nFpKsMJ6sInJO/d
ZrJqKz4z5kkhzn7I72vjy7AHmqju2wz3OViSthb5cpHpJ6T32pz/VbF489aztpGJ
BYi4qhu6Qi7xcBUgsTkd1i89+sio+rcAUYPHCXPwGTLkPOg5ohfFyLpeg2d0AyEc
j+Lzb/mj8/3+brIlPlEZxbWRHUUS9eJ1Wl1ngOr0/WEf1u5bS4VRZD1ZacQ++ksf
1IcHYYqcz6fSDUC8A/lcl+GnUVswgg4YXzfKxJOquig8b9XO5DMljJ+Ss5UbIoUL
FAobKo7LhNzlHtVi7QYzD5TSJMxhf6PBxa3lzThbW0B7Z45J2IEovu8YdkLvRig9
a1d+paFc/DnbiE2oWmvBvLTz7tJXTSYVuDJtMUziCUVOQS4aiiOgSbjXYRBBwXN2
sKaueiygJFPTOt6z4/aCn2hpaEASMQNV+2CVpTUgGmzUfkt6Nlcd1dznQWP13a/C
19bY7eYUgyzeJea2XxLK4+PuLnvWHo9l5Rz+1mnOiL0nS95pCwP2ZeTnUcdr+Ocx
MnxTNP6wnNhJd59uYEaTjVHD3I9ArPmZOhaH9/XgLt2lU9QGfqYrlqXfofskQ+AY
fMGbGz5bmoNSKXimtpwj46uuzGgS/lX47ekuHm3+O/TNoo+YExzB/wQgPE3Ez+Hf
TAWNP8O+JZ6TwtzCk5DlnsCXvr8+mn12EUWC+QFn5GvbD5zovf0UhPx7TJevED09
5RXfxU8XCY9tPZu6WjocWOmeuPTafjIu5qpyT1Qlm1B52laE+YcCBM20RLpV39yC
uj4WKGuUsx7u0wSmJbB+Qch7pdoElBs65Dt7svIxJ3j0UZwLatyKelAQ7K3OppIa
9TVYNCH2lKBqfyGP2Szr/aYMMhY0M0bcNt6EFqXmgbPGJ0zH5hbvEfIQGffz4H9j
VtMjNdA1pOiv7bU2dng/Y0II8rs/kHA0zq2uRBJw+Tx3BHJWNyDYLzliEvLapYTs
kvVKxWcZIsh9ct30vozlcXKne0WB/6T+L0kVgyR00zTGGRgnDQIng+tem24PBPcS
x/lDqgk27yeQ1QiyH8vV8uFur+AAmr6HiLcTcU6uKm5vuajuy//5M1rpMGC1AAHl
q8EmN9j7aX8rL0utGg0DkydVu+EJJChDWCpOywGvnsI7hMLJofe85v3lEQydvhr3
YFpyjVSj3MZamTw+P4n6SJV3tV5uSHWBDMppIThOX5KCL4g3CMDdwb5uxnjU3yA+
/CKPfpvrqxCf1XqxAuVXvQn8K95yMJXmTwouzOV/cVvhpXiAemfJQk2D78MHeq93
3T1HZ3Bmic7/Te9AFatiOcw2bIlHwWKTAxgPcl5ca30DDBYB3VdsZmfNIHHjOokR
dRyCpvt/rJyVrWEAyUSyL0XuB/2inQ8tknl6XQwHBEIIwFcSEe9R4WYE7YdDKYUZ
qztmcUdWDGbE193XcOmjFcTGHkVi+XHipAOeKjZOTHhA7jz1ynqMSGSFwIMUku6Q
TVn4ucGbBfwC6O9tUwwZymaLxxRkwrUFLK0X2aiOODxbVF2Qw5sqoJ0943eFqeMz
uLsG8xbhbsHetEfVFXtPei3nMol3XdFh6HfIqmgo9cVm3gpSdZzA5Xza2DoGgsZ1
1VOT9CiIU8D/+FlU+HlHfE3BnoAIkq+UiDHSRil2s3EKYOnj90BF7if0+hnNUN/Y
oH7IdLS2+yVUteJPsiTCA1d/aum3BPcebEH6z0xADpe/3TD5QoyrHDrAtw6Z74ak
xaZIiwoKNffmDwHtnQe9kEBk5okdCWTRv8s36ADijA9g1JqkQMs5NxEDCj8mdYUp
oJtfIj7s5t2OlkkSRdYbOphWutcMKCAoMA6pGyylG8VvGufrvC2dil6iKFhQUuck
jtAQL2zljWXvC8K3efmyNARRUCa3cnoXljlPetYkdB8wWOzimBVkiYtR2KLbMKZb
Zn3VcSx7MdN8BpYcCoTDFqzsh1XorxhaG57WAg1YWhgeeVA7bN8Ar4r1K7gxEEAD
htirlfTXrx7vhKtjJoFJOgRvO1/RYRbcHjjspuxufpLKn+xt4LJY0jPNeNRPEWCF
hnAa5mljcAljRslsApGd/ZNZmhCi1TvzMhq9S5/1de5VSAApz1Tg7SawLeD7cNp8
2dTE3qkodJN+UXv7z3YJcuerz3JP/u0mSaVQjBNl43n+8CDjUrT1IaoDVpcfQMiw
mjNDNTje6NscJBYx52X9JeGGfdOh/3WXfMDXhl126Zuo9/Zb7sTvO8M18Vv2VWgU
3ujZsF/NqxWqkXXwgzBUblj+82CoSUQwH1Q35VFZC2SNzBasEnMI7r+TOJMK6iIA
hbEI+FH6FyNsghs6pY5Zpkyxufp3sUn3ME0t+YVevObAO74Fhb/bf+uskiuWgWJc
VOl3xUp7Wlc0q380+LQcf0/6Q5NqfDdMghAZEYosISyGLL5Jj9GJduhLdHeWm/6I
9Ngcwvgm43FTfFbGSvHZaY2EMCDTEDzGQKPjSSzszMrAcysPwjL+55hdnLEpx2aV
I/R1DYSWljW9WW4nP8lRpktYKK/vEHlvfvlmrZdM2CIHfkrDjN8KCAJrdQYMk8Io
Mlyx34MYouoqW/YMoexplDYBlOatkAyYh83BZyuH9rZiCCMl0sayV/5HvxzB0dlt
6G3DDagyxk8ealFKc4YqcWBfsiEa8/c3GnsSrg0+/0Mqg9cjo3DU2dhYwQMyI2XC
afMPA6e6BouONj7o/zYb0dNXvJKnQP4HWFcV22U4PupLtC80lV2gUCD72jGA7STl
sdwL9Q/3WZiH3hNl5JWXoDSHFsnNzcbZeSjzZFQsG8VNVb/Ns8HqfueQoViGLodj
ZT/ejYFtysOzJS3G3/QGuA3KPYG96xf0AfKVJ+c0pryJHZawhuAmtr2DyqSPW6eW
nKYjNJkOUpXAT/8QEzK/br9wFzvOOVWkNcIrDCLBC0n1PFX/A+rLi7VdKsSHXxYw
YcY3lp7EnPApigdrbUd/t7DJHF2KXoTlXsrS6m9/EaBlL0wSNJsmWb9EurbMsfsm
MscBcioZaaIV+ATlN1Jp4cAwak+m4y/JOkIQUno+E/kvkWehaoi8bd+G4g934pdP
QZx28BcBzO7yQqm1yxVlfOGr9sKHjlukX4vcdIxuoVtpBNLNK7hz6NBYQHH9al2C
y3me1lCzHmfCil9iHPsXCFW5fhxreBFYVKAgDuh9qO7gtQtC6+HeVwG2VrSGw07r
B51TJ/q5uQPYRKKMO0RUnJFCde/jmcs8hMKefgV3ZEzsC9iHZEo3TXHdgODPqPtp
ulXfbFGTlkqa4OoTIjZFFHCbNVNuEaEpS/LvOeccmML0EsUe+f6U+n4+kTw6BZ+e
tN5IbeGN8gzJGeKlolb/IGN5VxLwFVjVKoXvrj1xtN9UUM8uaGlrJ9FF+ndFMJ9K
g1YvVoTXpTnexTNMczrHdcRMex3AymnkEltbjmGkHMusfMTUnX7WWnYMHeEKpeVB
FXNk1GwA9aTaBwdFTTnQ4EzipCelf4zofUXvkMLzoV4x0/PQHHgUbPeIhbCy7yYN
XFdUiPRRScNS5Lbb7qvJrT1RlQ/GwSUsf/H2/YVItwcUgwLIErAkDaeN7Wn30Bux
1lPwbavIvgubhbAqWqv3koWK922Xoug6Dxt64cfleB1a/ZyKt+hOQA3qcGanNstK
U7Cbqn3TbMZGZ2R0HYp/XDD2qQ2KeBo8vA2xPtMqbKl3jdLHN17979FokQO6VIUs
d9cxNjl5Om+ruCamJfAqCUjyM8//i1yLtgWkQu8gYNyXC5zV5MoZGLD7jbJuYx2M
zsU4CL9HUeF0MH6s0QgrRTza2cNaLY2a995SE6BIrrfNGG1/ECLQhWj9PdpeZEk4
WVdD8ZMKuVGNZYEkqfJK/TrF+Xb/T5f9e6AHjFywIgCxkBYS9BE2Fm0ohcls/vtL
q8KWmn/bZz6Z05rZujopW+vT7YRdOc+Sv6AutJB4lJxXOX8BJQxSBxo6PH+t2B2d
k2vN8qQ0UoW3H0FEoqoaUdXa+7yd6g/I88lD02Wa6sGTCCu0yLq6DR+3XO4OItIO
98UUiYUJU4uydzji3MtK6E/urPw8zFMeraMlj1McyoK/ZL/wgbafBei0mZZeKv4C
ELmCsqFB1XN6Fr8wMbw5KvKgsfL6UortswrlniMNg2CcCd6sgnJ8h5mhrrZtDpI3
QsVi02ZtimtJ4QhhxrToI4h12B67NtPtFJIjPTnVEZVVQtYRU1WQiFoMuH0NC+3j
GfIKYUoMuZoA0/mLunP8qGThmuM3f6iuwghPyrBnYMO2BAGrm7y9rm+44pf+mu6k
OiflPHD4Nt4Pds5PmK2r6WLxxfsDQYXwNz7ww0e4s0oV/l7AW/SxH62v0xvpYaYW
AmWsNaxiUOK2gsfXL4nq1hTLzOHifz37H3oNvHRP2BWM3LiTlimF3XKeAjaD2R38
i253JJ95Z6ZnSljoe5pi0S2c/W3h63BVXyaoeyLkGYA/ceXrwwcbwzXimaCcVhcP
9coR9me+tpNLUMEM3Z+eZ3KmcinprNR8E0jYXGeNMLOkFk0F2AHXAdiUL+VEIf0e
SHsxLsHCwhfSv3inLXY3Lz+9xAqVXN48VVIdPIk+F9lT7a+4erTVVp68WH3McWed
emtALBMZZHN+2Fyycnrq12r01tXOGSjkNDFqaytR8ujJLoTlLwmrpugEcQqcJ0aX
7gHSrkrTil3x19oAyQrV6pNOM7HkREx/5JFj9anyNIKtkrYXheFVboBclmRTc373
WuUFKKBpmBXfjdzzMdR3d0OULuJ2t2P/4dXCeg+DjSVsiPN5pjv5bRrDWrs2UjKM
+Hp6uchCfnhRQK2B41nXGi93aLWEoRzhPKcP3rmqyvB8B5p/sTkhmIsTWXcr8AYJ
7PTHFSS3c/hqm4B0YG/t9j26b5zoRrsLWakc9Q1ifHCfVjs3h4uXydefUtLzz1wr
25Grrcd6W41EG7MzJL5qEYbpRqoIgAGwJQSJgHrU3iFIajSyGvl2ilzGYDhF7uSy
X7WAxWX41s4FEhV0Ov7HtwYddwXtx2v121kK5ODU0MQufjjyFhCSQu62AXY9uvfU
ur7A5g9oWcAdH5Mw5ipn2jSMQZ355rY6KiZSjOcAabewPmoVvk61Nb+Nqnt2CNN8
rcrhTGAKZCLf9QVkvD1Iaqz/T39T+a7I1CcRviLZBHuqVidI8haDqoUsONXLJHPS
lLCAbjP+PbpP7P1fc5QK0StqJMj+DsqX+Ox8Z/Q1t0s0Ofgb9YldLLNc8CkjlK/l
6PMSms20L/OffqUVOh073M2LoG95Wjyg90G59xPQqKwTKWcKax1F4wm2mRhUTNxS
ZpESKRQjPNbXNU7iX32VNt+ZiMzLW96XRSdsm5dUW/CbpBEUSR3LVZvuynmkgiKd
JJ1GU4dP/ozndfuDAoZhAgIBKnZsGdzgfymQwf8viPGoJWGrHJS+EZbrRjt5UzYb
nQcfjYN0snEx1sPC1OwSz42yu70hoYzasJFJjoJhUsmjgyZaWF79lkQJNzrmeeZQ
Q2RZscuFRxlpNQDvUEJOP91Fk+i5aQ/IirlR3YuzGyI4rXjlVwDj20z1W2o5ppfX
i0V96p+y3aUCvBxAiTCtDWuF2Pb6w28Yj7MaG85WD0fkProCCT5PHy0HsBtv7XCM
1wWCpgFxbIC7xC/lm/x2JatZVgjUhYYX8KrumZFURIMG9i+lnrIAMzFmWmUYgllm
CTIODCA41j6eN+nIIv8NS4RDHkMBnUMRb/sbv4nsc6fr4283ePkZsFDGI0fEeWWH
XulYmAZ+mxI37QmPK26S6DWmcaKbyO3LOPK+XLEk3et3MZfRamF3zWdqhWZu8TTp
ZWk3tN3ThI05/uXhr8AYSumkfJLRWcW94UD8YKI0cbFhN3K/5TdDBZPNLqulDljZ
pWZ2YxhjQT36CHh5tCWgaAYCs2zXQps4iWYvPohzx3W1AZBIGaVAuuoObRf4wOpD
7Tp+c/zNYjD4meUDv5iBeNi98hB3VwR5LtOZMstBN9xkcO7YoAjYD/lwlC1IZOwr
rO8NfedxMYqTSdHCRplHI/i7ZLjl4X2BBAVmDDR8hnT+AYupJhqlAaC3jkC5cHwO
fkrZBx6kPhOgStpZqsMQmzS4jhotUt4o7DotHTlMaDg/E/l5MtqK1QaDol0IoF43
hHlNoqDEBw1QpwgBzzLumkIZNXJNvbJKGOcyuKWIL3I/6+lo1lqKzR4DMBJZ6vJS
Z0Tm19tOIsFL5rCuE1vkj3l6SOlu5ivw8heSv9PzFTJMF4UnQsqFRva7/yDiMmIY
GqOqMz8PLrCA33cyfJgTYT1NSUUAYa91box1o27Ewvub5JkBC9eXVSjuRtY0V1mW
nT06k8OWCl0QNZnu3KzEnNwlJUCvl1Y9MqRvJtvJ7BmqmIHi9zzA4PrsMvBlZEqk
Y7yT99xInRKicZMjkTnfC/i3mmocQ1OCB0h90pu35z4tCCBOXNf0j4cgCNwCgZS8
ZJwmtCrAsI3/0Y58ZLqQkSe6YTJlH1Wnb90tiv8sBWXRjjhp6wUKafPYFC32qSad
QQxWtEZ22CO4zFZtmmjY0ohNpMQkX2fyx0Rdg5m6Au77lGhTm2N0gtmPRY+NqqeB
1qniGWaw0lKCb7ryE0mObhbIl/CMvJf6Qv2VakXx89RzxiREzpe+S5nl6UGVawEc
Lg/Gn/ZcYs0+dnNmuLuVmGrrDV2x/qvO2Ub7Ve8raoNFzstQ2g8Y0sZMvGg7XkfI
7QpyNbj9LqC5ytMsLnKemt5MgClmQ/1cTR+2Hzd/D1b8N4aJD9UF/tJQktvRpP5z
7BSNo6HZO4S89pIF4Y8MAHgIWzTd53dNLw3C0aGFfGasHS0iUj8+aLMTOlfoYwld
vyWWra2XxNlkNESxHrIsoxSqlJbl9bEOT/0pAtDaXGZlQggmkcEDW9yYt1ydmkrE
q2o9n6NCNdoIkrGT7PhLciCzAIEYrM9bT01YaDWuZ2qvXbb7wfBMhyQTXN+dFTiQ
MI65HfmjIisuofoiR7m8nGi1CoqqENGl96lhLgdP3b4mT79Ba+tzE+MXFAMj7kdI
dbLnDSLLCRtmq4gGX4ETgUmXkZq+oekZXecmmvBDBrSC+9X+h63aaFoxki836taR
L2vyGhXT7DsdNgNfmmyt3YczOPGHmh438OtUhNWN2fmGSELOcaxcQ37oxPzNAsNL
ydCOQ091FWtDuujqWBxbgZd4djJQ4H14LC+vCnI1yvXm3vkjg9ofT+coBzflBfzc
S8VcBh6Eic7LM8Xk9m2Lm7cmRj6xlb2xsNhGATEiuyRZpexcaiwhmirSn323bruU
abk48/Sf4LuRoDiB9bWJ7yXDKZW9qcG0ooJ/pKo27b5SxSmga4HTbaoCunmmzhO/
tGnEbONTySLgdTVI/LIImseynn/c6bIN5Envh1azOYYe3evoHNEoqT6XK8tbiDiC
0OwOqjuENMgi7h5X8JPTjwc0mWrJAcz2sgIm/ZRzfGVVxTWDFLBmHPh5aGQH9w2U
/xj9ZYXgTCoW+ksV9RYetIXQRhVWbCGQZ5hSDJsAK4pUgKE1veMCXCNy5S6gcezD
DglODY3LdR9fW+xZ99VDc0b0bThCQeayM9rD6427WjWp86mXfoXnaeI41f24qnK1
dkDpFZPodlq8yP/nUugj73g7CQkosQ7pGfRz2DC0iukqpzSn96xor5C3i9YM37/f
ijqhwSaGPvdcfGvua86sNXiagU8C4hyZ+RKVQEEOGW5kLtbcrLDtNyzn4ltPGVNV
2TRmtpQ+7ZVNOd3vMCV38yILW8ljWgE88amhp4h1F6rGfzicDBopAipBmNNWZrDE
Mf/cJfIUCGuDk1czsFaWXBD8LCqMGJhWN/NFXEZDvd5t/LSVMjuHZa9UafNsRRjg
CuH3fExct4/QH1zNd8K6IS9Y1303pkcYG7ceCqlpsrv13GYievhkBJLieX9qWQI1
4m2VnJmIq0NUTGE/vn289NWu5nikpF2IR0ytGBMshgMkbiIbWaUXaLCQPfpZ4bJ+
Ep1TDuz45jZeqqLgwdnABRkj7xAYtn4p9PvnPWcnI4hd2jvJ9mUmmp+ejzE8L1tg
fK7C00fXU3pDyz/0Lota4EWX9g++ZnM9dVqnCPy10/vy6Npi71bggLH0Sc3Ozp+B
6niGG/pvoqF3t7R1Q/6f/+sIPFZvYqy9HLVUiC6Q1N9mYj384rCqpy9fFLBgvxhO
Ze1NJKBlJi93xjQPcNbOC3WDYmUfjJPxufmZ7GC+B27bF1xLWvROF1qb2VFppLQh
mscFlnPJFHcZi8vvbvRO1mYvXxj8w3tnAhgGiR03/GEkOaNYDsDmccB80kqb6YTC
DNhhVoBK6YIvwXvPAbEtk+6SKOYxjr+j4Dh4RSyRirk4NJ8+zH4eyWzvU6bqx8fH
7C1D7lIShlDjQRYYz8K65+d4sBbz8BaE/ohVS2JP8BRpJ+enFJJMv8ldOnMMx6ZY
2vYNeJkRZ8JnPM7CTvlrh4DKR3oWRfygESGCh2quEzfx9srC0bis+7wUMFFLsggT
Un57nsp3c8GJBq1xgwvHFbiQf94mXIKbEFIP7GDzD8XO3eNOJw3JFEM02MH7epM7
SOkrKEGV4aQwbux4DNXbvmi6Up1PE45IfFV0bRxwplWwiQ3Tp70u4ejt6UAg38ko
DxCkLOg7ndXMmXC8iUGfqslJmqzTZ5jhqraxJ30oz/naIgAxLI1NMhIjIEjDaaQU
qwEC+lvx5z/8hFZqdufE8BLWglLUMWHAt3sOBzEHDczxvi1d7ciX4ZZowR8B7ex+
QOOOUxRb8Rkoyo3AeKtH5AWoFIxgGgdlOG7pqV3URbMI4bzlkgFporqgXh4b7pJk
A3ULInT5X1eMIEHkZ7f7siKB3qYJP92/sh1OTsouwfFO0wtgOGPIEnvPYGrQr+sQ
8m3dnN8pRt5o7mroYjt/8VqoT2nRvweyKsPLEi+kObKR8yNkfFv3M9/f5dyEOGYe
BGDU/EZsxWiFFmOmGgjx370NOTuBO2gkSMH1TFz8/Ai2Xo3aT/SapQ1c/s3H4C4E
iWOsRlVly7s+PvVmvUeojXtgFL8MF3vmGGhYwlNdkGPMQFRMqomkESArAPcx4qud
fA2s6BBrSX3JkVDsFnHu8kCuQdtWQpHNz/Ec/EvYppDiOaYqThU3M+IEV81Ep/XW
FG9dtkD4SPng51v42i7wlELewZIJArSu8AVmAttGED/0jw8eQLMmW93eQpFeQn84
8vKao2dreV7Fq55SjgaywAkmhKb99F7MZAblrOzgVnUeaLIIPL0qm2uNRhq0HG5h
nDFlQ7j8cOZzrWsXJB2D6A1Axt8OdwgDRvMa88F8i7FBP4Q2PC73zpG2McVe2KEi
/Pk1b62yz0uCZmF9LXYGcndoo+nLjNzZMub+0/CTSRDIou8g6yFbKn1crTzpHE+R
kY1RQ7B8Q3aIaIYdkidtEHwB0N/Tnj1ZTLcvOClEXcU63zittmHzmoWSB1/Ydmvb
SNhsBdezmvBxYFJXIVzy+VlMQmBxpDPEebOHCVGY2lnexb3bRA38MtXGLdZcIIiO
OiNHVAI2TCglk9PHHuzcUB4OLupB4qkaWVTVPGgKfclye1V4l9ZzCeQ5Avpy/yQ1
rZZBubXke5mx5z97nGBMn/6O3oBM4JiyOUGfSo5vWxuqGO6kZLnGcbQbNVipIBtf
KYR635DIh5WBQNYHGAYxv0aSTdsmhkePA6n53EmG6RCsKOUaxQjpoLj/pwnaZUZf
2T3lswWu/A9xnXbbXeGTc4HrhNf8tF+8FNOZE9IUAm5IbX2BkLDdZhs7+yjG7DAs
euX8E1CS+ia1opAyKL2KJbDGx6RHej+IvhELk9UsW8/QCSvBR3lERjje1gDZO0+6
cmsj4GPd3RpowgRN66VMbwAZU41hiY+04TgTAUBCOVYG0wT5YWh4bXm1Yu98kN98
47LHTyYXwHIHsKMKtY1oNc6l1RB3VoaOsbLV/ALxKgoCJwW5DHmY5SBw6EcrL/Xy
O0RxrZ5bui9ar5CHgPTzOoKGOpUTUiRRoW4I/mwhIExgCRSx7yn8CRSUEandcLmt
HHCSO+IpT5GPeuF3yvmBoTH4uO1P4IuMXfEs8aSyJdpjd4P1cJhwtYorplPTCQ/i
Lh89CCCcrvTcr4IGt1U09mrGV/qjxBzuvCuF4Z42dPew4bEBh4biAk23GPzM0oeL
ZTaGetgY+6RlwRAoG+UqWgyYk7tlQH92EyWhOx//WXGpHLaSee/4f0HgQtkNSQzb
PWfQPnsn+swM717Rv/W0yIl77L9zZWl/H91KaIZmvyGdbwFwKYg3JtIBB7pXiPdb
mg6p2UAY41bQMqS+GAQ+YroN04gstM+XPyFXM++NieBSfGlbNUxLI9UzZeHLjIIO
UhqwlMrNVEdu/8nSAR+hwzDiljySkUHa8nk5DrA7h1L3ch8Kj3UzQ9XZbRzcQkM3
hiiuPsZxBoF8gIhjpxu+wfXug7tUI1NU1/+FEvv1gSfWNYt/siDYsbQIqYB9XAAV
Jqu6Qp9B4Sh1VcrLLAJJB8c9MGtED61VRFcT9rFivF8x+pbOES6XEQljdEN6YUH7
BYvjz231QDFOu1Pd++IYG2HM6yYwcPM14/iH2LwiaSGUrRQY/8ZZCv0E63mH7+Xw
cdOU6zu7wM8hLj0rBncnX1uSkgSX0HpMB/Nwv8S4oDTHnUvicMFUe2UhNEQPifhr
RK6dnH/fCeTOy5eyyfNdVGUq9wOYeEKLQ+8J4dBplXGEId6rgY0uPh62+c2YKRHw
wfGhqrt4kc3ly+chm/v0iAyvqgWNEej4jIsElSjCnb/Nd/UB5IURVAY5lf2HhkyR
rt8XZ1PFZXuYEgJHM708hV+guH56oCht8Ic3qoDk3g/Cne8G4cTPir4yAwPnGvoE
qazuKABggPaafpyJDOS20aJCz0Ggo4epQ1a2/jZ39TWGY/ZnjZ4RS+5Iti1zZVRY
F20F6toN9JcG+89sXAZg6g==
`pragma protect end_protected
