// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:52 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
qkfNFpT36wH6nHGdWMpKKbhK2xtYG+1RHtMmE9kFd1cYqyrJlGK7LLbs6WA74sjv
LV7kD+xlTcj2Io+stjF7mXBB26QhPJfpqJYRaHEbradcofHeBWPm+VEFQyPZY7aC
GzSN9ULv9pn2uzWm4X2Jg3RJWriVlTRL99aTnS4mRfg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5952)
+M4daXhm77gr0fUJEZvdDxGGofhRzzMenavyvMryzR88JdUO5/R/SJ5+5A7qXZIx
K95lesU4FMtlZRBorOn7F/tStj2voIL+9sISOZG8mmQtYxeXt4zPINnEnEitCowS
MKggF6GbDLmiQBnZcLjVDdiHq60mnc9ZN3f/T3H+Do52EoX3Vmsr0ZclPuvJcMFn
LBINZJ0nzhUVo24TkE9s0OoVC6aMNtTebhEzD+B29DDjpLrarhLlQBuGTtAY+SdQ
00fcAhln2R8VBcHu7E+pLwfaOYRE6RwKrmac4OOQMCkhntm7NI0xoHoYVV/ch8ta
ouoqBTXpDLG+ft6Bb4MNb725wSW1XGPD1EiXeukwEsfrB3XpzHs9qUyobqKJ0NrY
xj427a4+x6CjBgc7synWzJY7iV5Re0W+1LY0F5Hm1i/PzE9Iekgmh6AP4CTp7KH0
ZIKGoYX6ytpyd+AV5fzIhxmKB1c26V5T96u57hkvW1ZcaTVLL/UTlz50SfGNiCpP
nsR4+vKuLKvSCMYPpdM4ZBa++KWeKTdRXP6Kq8k8VcIg3ze5NrODrostxHFQ8euG
GiD5CZwJaO4AjIczRzMN57+yZxFxopKkFoArhjrBj8sO3zIkVNu8BXJo96U+pli6
D80eYiwAe+ykrSnGyv8QDGJQPcAXc5I+MXN+1Q7Ikn7a/9qV15l7ZHfNIth+Sv35
7Z3vX0h5MhucnPfQrmZuGwxw0LSRyK2xcv/+oiYYGiWqYawp6C4ZWifS8ojqEFz7
o4ZRIx80fxW/N6tAm5O6Rsa2UE85nFwPWSX6MRCzFM/Hi4cv45svdhqnsRQb5JRg
GO/xhJ1ZCqT883oEAhQsP8U74qQ/UvM+9JWaNEki80nQpQCTcpzWyJjfRVVeYdK0
YV9E87l9xX4XxSexs1qpTlBnA5Xha8j1gM8IzuMe6BVijFEwMhBG5mPHLPUB5Jmd
DSmPC855X+UGuZItWoXuAfrbGL4EFiPQUEoRoVSzp6XhF83PjqwUYecxhGgwbW76
4XGF4dR8eNGe5bIfdRnRS2nssFVzQJgWKW0mhVhhxsW+VdFsNI41EoWGAlPCPqmE
CjLOrjQt6FBnBcxn1mgDJFPfpXsPJkEDr1IefvdbZ+10ujrfPrvZML75Z9RzXqI4
WwPTDkOrXhFh7xRxBvdGpV+nWIbEeeezDC1+Zuvj6H69/MQed4aEng4vXlWMHhBi
o26cs6KBnp8R+2Qrk12Ot2+igT7XuN0XBvXqIUYiH0ngQXlsv7TB6VSieImWrCuY
rGelAQefwYgzGNoL7tLpPUGteH96Qsd+9xz/RvEwtNhhen6T8/HLdeD0fJgwUTds
/VUcvAC9avGBdpedl95ezOXWGsV3ZkjLsYbJfwjQF6FK1pimJEXyHfvIGdxoh0q1
O3I+m4eW92gHm4Yg/l2hLfeZdvKOrrcPPXl47JWSYXZf5O38YYU5J3FDmF7W/lhR
lbMcqS5futGHHS5QqLGrCMoFCIl59A07L3Y07GMsXXFkfWdkbg93G/lhCgKH8jMZ
Y5QZtwHXzysKLa0J7oj75oOQwuMMBqcJ2a2JlxwoTlifOFNlQdLMEV2Gbyjhc3ha
4dbSr4InMkEyXrp7Fx10hntKQsAb4MaT+l/cQYxDiD620cGrHOgZD8xcXJax+fEi
vUft+5iV+fm8Uqst636AZkBUEqFjbCAREbS2JkWKOJJUee2I1kkqlfkecaGyCjCq
Vf7Rt7VlUI6RS0Hj1l7oiYiMTB3OJwlw8Y14+tUOkOUkYW7/ntQr0ZqEIdc69tf3
XKpjfvQC1nJy3svjPKFEoZbd8TgmJ8mXrwZTVdmC63ODmsVfzumWaNTP58uUkMxW
zZgb1wUUONqBuMulNff80knhE7dcQa1bSY5TNST0yihyJ2OWT4ab6W9Lcs10ioyc
flnXSdPVXPqrzW4zrDh368lMxziNPmToCP7Ey05xjKagwloBJnSSKpPwuhVCmVr6
LPKBdpp2xtOmSk9l7vT5zaAYE0uEtM+KF1ddE/2HaCxB6SL/IE1sy0Zh5ybPCqYn
Loz/uZi+w37/60OwN7uGCMkTBipxhlmX1zGBh6TLgponMq13IcqgqRDY+DsvOHYa
WDak1zn8J0HrpZPXULJtBouVWId5LAfruiBNbRHTKpPbSA7wUGH23i/qDk/8zRYa
sPRtxJil2467oklKXhzZdpntRPWvfpHWHh6Z3TRYD7kAkXfnt1qWrvMITok9QiS2
A9ZVeHBxxIuhKCA2eJcpGZ+ETH5NudjJhognVY7O1YcoyExbBPvRdIQIzCRKWeaq
Pa1Qa6Nn3CDPX9ifjlAlh8mey4OMgpwZeOueV61ksiyZPvk7cIez2F3Ggmt6MJcP
2Zn9wbEGCh36ZyfjSBzUZDXCjZPgygv/tNz52Y6p8NdhuhwKAHFnRpb8UjnK94HD
NEIeVHWhlNfm3+AtE2MRpGk4jSniG23uKJeelebJcwCEnWdqXICHWaG5TxCt3xP2
GuqKVklro0uD6rcbXmL6VVbh3bDwnH4jg0M5p2JkYbbRxf7az2A4fj/ETA4VWX1R
kph12gOjYoKkOiIq4apjNzKnVRY6U5Nn0l2Hjl+XYycwdaC3XvJCjjTPmotuA9PC
ccCMHzIH1/j1k8qRr7DztGYvcTvoNxluXxgHICnQwQOg3BHXGEsG6k0qkz13zy0j
u3RvwLRPvWM+oDTnQZ3HQ8eYo6s8CqlfXgMtxPJSkmFPhe++z+ftMxhtaLkHPCeZ
TAaAYQUoBQYiLBCb1SBlB7UjleyVTwvT0VSS6H7SZVlGGRMbj+K82DlKgS8NdSDA
0NXCWJHd7fanva0S7hbwBTmfW8dO14F5rJZapYBjpVL2y2T5TEcJz0HwDIOJVIM5
HXKO/f8ShbuVGS7OVLk4xzn9XnJeugEsAjdcd0EGvtgw3PB8iATRIq2aDE9Rfdg9
vABTI4N7I2Bs9eVG+yuzdANcxRWyQ8loW3OfQS6y36xElZk8fny8yzYa8rGATZEV
BoJjWvB+3HDGRTVF73kY8uq22UCj+FyXau5bs+D1diCsUKdGYBG3Ka2DX4ToA1AW
GR2rAov6TbcBtjU9zkb1R4eSC14MqmUAYeN0ZlEVt9aMyViz8EtiIL5UAH1q3p3w
VI/PJGp6gxwXWKAO0G5FYJ42hWnpcivp3v1bHq6o2zXWZBGipXc4rhHO+Ez5ouar
YsfSp85pXSlaZz4dSxYatTgqfKFE4XbY6DjW5Zkjnxirr0STbZHrgUprbFD2hehz
mU/D1t3O/TmO9/Yp7KF8rsyi4LHr+LPejM+wUMg2+pgi4C/iSc2fndDm4KV0L693
pXxLaZ5ebUZ9dABUA0+x4sYYWdnaCY8HGLjOF8uBIEyIsYVY2mu4POd38audIO62
+n4EdrvYuVdkY3aWjRauOH2RgrebbY4ProXcnDPsmZXR5DtMxB2wpPWplmWt5WWr
Vy3RzkUnFdyH8GlkkVCXdZki+WDWFJgrR0aCOXarNRJQRvfuN5Lf1nrJlZlBxrHC
5l74Uuz1JMY89fCxv+pIPfDtLPT12Jz/y2gU57RVaPAw/YpEsrn2M/mNpnRAgnjb
FyjvM2eNYk6FWXNhc7MLBcnMdfq3g/FIsTZybIfE1hkQinqS83Oq+ikr829pGft9
c1QnnvYHYDjHmUo9/Rf8zChh7IRwBryimPF37Qqdpj4oyWQqNGmFr1iNfhabwFZt
ayxt5tu0KeGlDFFBgO0XxNATFq0wdIEx4RI/qyBa590kHCfBOd+covPO6Iyk+Gg3
IRfbLerXTwntJwgy7fusDMXlz9SCydhf742BZnncOz0hYmBOIaFKwNgBkN/d3Jbv
1YQAjlT7aFvgS5DqAdFk6xyUpAog/x8klXWt4SStCLiuA0AQN/Nd8Btxsjj9SmTW
wf1kGUklETe1xz8dSKZ979T5N4ttnWq6/5K5nHVVEDks+Oc/IZNjcBy209FbG755
D5/x/wErQhpM9jpaQq1oiuMJHcJt39II1yN7F+qXBaSM8yL55s4wEozkNw8BeWyg
NbOrh5UhWyNwU9a5kZWm4IuZCzu3lhtMrdJfyenilH/KYjEYl8M7sEHa7Cq2PTYB
DjKn2WZnkncOYWu2qZLl3VVnzCip/YQ2tBgnh01SU8SWyhsRj4LuQixZPVvOKCat
rfUbaSekokQc21UnWijQO2pllexZlg+vWVeGt8dFNHfhJb4220Uvolj3LcVPqTBw
nQgz8gJA3jWdvgA+aCph1+D+P3Dacxzd5pyTlBEdrPDXrpJiBYOqJU1t6BhXaoLh
/2GvnKfRWW6ENa16mZVkcolEwCu8ouL9aPHHWVwcnHg5SdpIss/RG04BLIq9DY9z
5tzXUH1qGZzBUwiHYmfF4fYwUAgwWuvD1hzAnC4Q9fTpLyH0h2YqxiS7tyVsjNUj
gRt3ha1ffhoVionHyRRUG3koOTRc7srh18m4EIXo2RBRzRjSRwWpgEdtTDi6HH5p
7PfmU4s/j96doR/IYQIqplDRjG1BYjjnHvwmzuVziqKujm2dEXSXyie8l93uc+k7
ssE3ck0GLMtqz6qdBnLwbkGda/AXp4ceSLSNx0A5r/A5vof/Aj/69migxygdl/IN
ETiZ3b6Oaw7gZMQY3YDV68noQvbV+L8ZLSiqACBlQh0Zva91NrqwPUFOYhAZIy1M
h2T00/kzCEZInaipNTSUipRx+dIFBDhNoxCuYaYrC0PAkHL4CzxlAyrCX3bUVlmR
ToaznYv5iDeGVCLRiybCSfft3MwCXxIKX3iRlpv8kTdfu7oaID1bh6/DQVAPfpn9
vKAnsnZPLWlfk6BwLtt/3DEQSPbNi7CEnvmOy5ghAWARrJmNezp1mnBGyDK9nTfu
P66g5wzIRmJwY7BoLfEv+rzF7fsrj5IW8dRkTeO9zRvQ+YigRUotuY4FFARCpgid
b25skAD9phh5ajpjNkgynEwDQcgtR87NvrG8Ts+TGzc+WxAEe7isemojdhlFmz8r
A3J32Mlxb7F30RyrQaHPgAxeHQpnv2HsWZJOV+/BbHlh4BnxHhAxaa5utrSXerYQ
Qnl/3TYxheopn8q/KV+LVjk9Ybg6V+7mjJnAb8ojHJjLyKYzoAdr40nceoFXYLxR
MOHKhpaLP6vEgoevgiyOiBkgqu0ROjARGxSRofpBEP9hKd3J/HGucXvcXS4CjP/D
z4JYzALp7IJweuQNmiW2SFopuR12EHLJ8+/HLLNQaMIy4biqQQLJz/GZPHIL7Lg3
RzhMVHSwIkGnD5kd+avtYK3DSUPaQ1JsNMfZZFIeftFehklpUNGkuQky5BE/QB41
oTqns78hjua7fEDAtkbWjTTmUo/cj6zDDmpkg9aeMt8wcGQGPlIE4L3FabwM4gyz
X+5TYG8zSLJdy2nwqBOoT4s2bD8jx6JpQysXg64M/LCS5y/18lnMJB7liVu40aTH
9puwqS1Z5o9/UnPJTnK2bP9cyg9uoks593AUbbAterQEaG+ICUOqYCNLO9PpeEtZ
yzm6CCfVRfrDk1Afvy5XApKk0r8F3oY/HqSr9mkokv+N7iCcYmVunZdJPy2Bzlty
Sg7WA1LcC8vtrpGK7JJNMhUZQwO2lr2LnD5ihViK4Bm4OrjCoIV8GYKVcxs3uZcb
HItlpkp740ovf61QiSDtT6gLRPR2yHubRnNVP2yWkGvPwbXFS2ZG/MSQkSnoHA+y
4OY3EF4fE9S2kUY5kIqHPz3CPtrvnfLDnxckYqCzjnftroNP+tvLkBaG9ly99Js7
gej/rRwVjEe+EYdDgNaGeD8jAvdtuW6l+tHBtlKU7NOrHo3l34UP8swGbmQQ+/jH
QkcQbwxcbC77SfrAfSAARflMD+tgHnzgytRDah5lGaB2v6jbt0JcvoYC91UbYqVZ
oIMxkF7l9F4CPmr3s7vZwXTLlomOKPvtwIYeOnzuI60CR6COwgDtX56vRtgtWC8I
D+aGxPTgJ1L80WTmGlRGxYT5yLA9Pgha+R3KifS0Vr8mpmN0536bgOmxhhl1kMx3
D/8rCVqIphbkNvJ1C/CrocSV8N9bQZd5R12KDOLz4aUaGUQj5LErpWZhlFHrrNBu
9XWzuuoAWlmr+rIPFLs3bwttEt2+ZT2GJxDP++z6B51A8RfbSGp7EIk1s4UnrVSO
KM/yZ+v1LWDpNnrPJ7sdUUmARhFuxC/yEwNIVTFKvT4mmMzMt6oBRUaHYhUmRoXx
Jp5ClgSk9y40jP6eWeHhFWqyePCCpqaoU1ztNIZZRADRLEGUtq5751oYHVKk41ZP
oJHdwsOwvlem3InhHn6IwsNKxyR45d28MIRUIYTf9yhDgcss9UdCWTxgCizRwGu4
Zg7dGpWQ8ev3ZVhn8pTRiIzaqZnkrhWc28J50Id5SrhLEM6O0Sy0o0CCcOB0DcIw
maSiPvnP9YiYkKa/vsvMrg3sgdfPZOmzJQc00DzqMKFa0HS8tlFUHD+5rjVBtlfv
kmz22FSp3Q7nFqW9tBqq/fxljviXV1u3fDC6LY/uiVux7fAY66a1Os/8fatnMC4H
Gp+r4nozlSV+BJT7+iq4iGRhwuFfcZJTnqs+F6BytNgjJb9zyXqipJD4OCcbobvZ
SKXZCTWI9T2B4Bfk+YOqSABB0n2mcKPc253o9EhW/UCmHodA9x97sllaVi8EW1gU
HdfiP8NqeryE6xhg9QSwwUoONhVXDk4Vf2t/HkCIZGfQSejbzoL/oMHggEbM2ZhH
GqAQP/zmw0ZmO4LRmq4Um18gtolhAhZGWWdsL8Hadhl2wT6quSjko9yNCNJukmh+
CUZOoSo8+2F3241/eUoII45TDW5Rrk0xW2p0245K4snits0hgwPjXxmwwDyIj/Vv
qHCqm4NA4a2Ashhxkulw0mij/bfM2xrP9f4Igu2cMYWAeB19raaoLVw1xVB5DgYa
xpILvKPshoeh3o+xyb+YBMpQu52f0J8xoYx/NplMaHphAdxZvY7dfpJT4fbcF1VW
8T8d68+Rjf8YFpsTPagF7zcWtcSMRkhSgNzwMHgU4SFm22alhDxLnpnCSBrCBIP0
4FJCxgkJP16aVgrOWdBuLMCdi5eMQUwsQUPOvRoLq1V8OsiI7KwwWRfyKJ5JIc1O
//xzkhXcc9E6U7yzBifjty8TlmrhBS94XfwIMLB01oD2aD+eHBIW+8LOF3HSMGrp
73hCm2y527H6GNo3AsrgS/pjJQqoDVjWSi+Qr96G7TZuUklP8qOisOGFkdt7fTrH
O+EBTqfRB3NP7wQ4wDdwIz9ozLK7nVs18caOMjFQ2VEh7JmNsOBwraf241N/5R9v
h0vlIRfeTer80MgJRkHcLHZp2y5B2knrog8ziWmekjOVGpwS3NkNlYV1bkW30AIn
c/LQCAlZEEGw2tjEe/k3pF+yusq+RRawsrw8YlMya3i5/0SFZfNEIadLao4WbADF
Exl5Ys9iTBQiryMlK1YeHdicLsa3GZYqmOHyfzr8s3XB4EBQTZl64LybaSl8dV4c
OUiUa3g6yF8R1E1iPk9kInxCNGb1QjP83bwnzww7Y+BH3r7N27Lv5Xw61qm4mZAY
u3zFfPBIyspCr7hhS8XW+i/Br8CUok9hHW7wLXVJaYQIZbSVxfhAvRNrqbD60k4c
hQzX12LU5Vh3plpyjEjuys42oJAj+cooxeX7upKp1DMr8g7zblbdP35aSToSCVJP
laDw13p5Pkz9qxAWvtbWUino38EGuRy7VUiNKLAwXG+2xTJ4lgnyJdSB+6oUBcSa
/wTSfSprWO9MoaptLLZ7Ey5sHfO3+0/JNqWIQf61LyDrRU+cje93eS6n9UaLZi3I
RCFsy/LHbvwQL8tm8dHMnx7yYj4qwAGZTdiIbxkEopgmM78ajvrORFwKwBERO26s
dBUJO7zeEEqI24O1GPDzYL+f9PyyV/OoidFo2qLnml1LgNTRsPHFF3c7C7ht33Uh
`pragma protect end_protected
