// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:52 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Q2aphjJgrI4+vIH26ddm+I74sryUTnkPARISTUifnZRs0yUMhbt5HvqTVu4C6Ecv
h0Lo6p7VyGF5J8Cis94SchrIa97oDTiUa2DvtlwYCB8g8Kw9wNOlqQLGIxb+RTIk
5mgYjhcXRzbRVsaq8pAh7RWLHG+L2eaUrkAEa3qo5RE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3216)
VQpIrUUmR/SOFWTC1kSTuBPiLtHqtHzM1FogtMzhMBfzrxBc3EL4JLpHzvCHoMTp
c4xltucB9cauyzzVF3AbWdwDhpXqKs+FUf3tM0/rMLNPZGUYjZFKzu640Kv/s/Yt
8Shm7b9Bz8O6fzunB93kDTk7NligpiFQkFsgUXvaYTJGJus7DaewUBbVP1dOkd5l
oarTvfl9i/PQQ+7VII09AOstL75SM6Ig74Z0lXsoFanJY4Mvtuur0jRFfN8adUPe
olQTbSpNhFw0kTlIrIcpWYcV0q6B58LbHMt4PFhhlwkps0vkONN/hDa/5VqhpNbl
xol5MyZ+ce5tNNJpRQXY+zYl0FJG8iPplVEVxLyv54i9DpDeyC9YCaraa6SyQ0LX
rEJAdbChlCzAQqa340IDaFBVYFgUuy59Gb5Q+IrHo/zzFioAYcksqgTc0ii1Tshm
nyc2mtYHYHqKhVrI//UKJszxhUrdVAM7rTTIBCUJOb3bo5lM1q2AZMCpGRDayfsM
rmEc3mb4V3vb4pRaamuFFfnnxfBRFdM+bT216pgnpNypZ4oziByAyYZ4N5o8eAys
ekH/ko2Pkc+iH9kvW8d5Z6qWIGIcH/+NNlfnhvHwWtJC3WWjk4uCcg518yr/IIOw
nLJvlNMLgaV4JSJLM9KKnkfOBmEZD1ZqhEHjeC24TWz+BCyLiteG1r4jbKn/l8Sd
m6IGJSbn9uI7NfqrtYVilWpihRtbV+SlXLSiOsAwL7QwiEG/xNinnX/uqCQC6jRg
hMP/Vqp5eLl3V4OX/jEOmMwy64iD3RSqZQBL9LYnO6mmONXE0LjP0QY8HZUkmcq8
W3kQ3E9rrSweAwDOOqR7vCZAGNeGIlWRQbpijIgn06X4NH7TWi2lVo6C52fQ12p/
XuN/oDdkJRoSfpmz5tBMU10r1FJM9+TLXKKdaKGtDEhy7ISil+caL4Uwhjlb5lxi
ez4+17uaardRnZ56qDDksScSakNdR9TT6pRaF0emgviWXfKFBNPVNm5xJaokkn5I
PNJJu1hG3mVYMfB/rBIWmnaiNyHWxe6ZWXJtNcXmFfuQ1bsnEhB7Nh0Q1R86IVut
6XJ+/X+htVB3Zg7iBq+l5iO2PvSpfBpwOSNDjeCZkkjM/nxKkpCx/Qbr6ezALbOr
iHWZMKe34lodM/X1g8wV/4aD3kZLut5YnI7z4YChbunXBHcId1FmI/pctwfIy66X
ldbDMWvJWTTGWLSWAHLozJPegdCL+4TZBvMlQrQvXyCxAEIquLjEx5AL3S3X5TXy
uUQcMyjmB6wbFzJJO+LITHiVEtlDjN7SdIgHUYRH+RHQ615rEnEHyfgQg6fST+zy
LXaVwSQkWzjgI5My61jrLSFlaVjjs1VtibpShxHd/XfWmlQF4Eal8yqqPbP5RgOP
xkmtNE68V1+QlfNUSD72iOT1gkPhaaMgzYUBaC6ByPOqcUO0KpP1AJpdKQJiCiPB
esdo2XLwQdjRZ4LWSWHRAV5gCR0jgBu7rJvtOWuDIfbQ8DjsPs3j815G/5KkzEb5
omkrqifN7qjsSP1akh0f9yn+ekYbJqCsx9n9Lnze4D+eknVSC66U8NzrzAibCdjb
DOLTteWqbYdamt26zn0N32gLHs728Pqdrg1e3pLZtB4BNCwhuxg2nKk3HBbA6fF9
LczArj9NwCZkDfRyikdzIHqgsEy8nr7kGCHd3MI9HN7wreJRPS20yIvilH+N2Jq+
1zbwgUWOyDMaF8XWcieHxrRRMGdbHRK9rf9em+lzxvSgXMFxUnpK0bi0YO8sxDqB
6wm6WP+eNSY3B0o9gndiiqszDMkvRaT8nPH6QJtfc63rIaHtgnIrByaVjbSWyIe+
wTDXSbus3Ige/FFIy3JpbR+yEGwHBDQqmlITJc/BeKlA6+uzRAxa4ryzJQzShkkz
ef8sY/uaHRXTTWYbx6cKOTsYKAd/pVOArLBW5KH+DRv44vOf5Wt13gS9ggiJXa3/
kqrUeozr/0hSncQYBwXvqnU10zOEI/CFNi8V2q6/Xtcg/NJT3hRA3co+GaXE5slt
6QZBsFJeXZKl49IhaaTFXjmeKZPr1SkS/5PEWBnAynNnRhmeOfagJGjBEtQ0afBC
lrp+PebAabrpD6NMyCeb0G04oxjI4YW/tpEcU7pT1Hi2lN0hmEzpE1NiU2J+OP0E
q0bZx0gLzqfT4+KbDD55usW5F9IJDEDQLVHabc37KqPGJIgIWJWvpI8dRlrsc5hD
JyCydsSNqnqx6CpS1lv7K379VfTKP9tgcXci/rO2xrEgO9xxxIbRx+aQHkulCiGs
IlpUHyJekD2RWMyqQqonTNKxvd+eCD7ruJ+bQ4L6VCck7CruIBY3j+tPJ09Z2LIQ
PLT4Cy6G8unponU1gakIjOikbZN+wKr7XYWbeZNuYhZLebM00ksJ0bXJw+hgUsEc
nL1j9g2t0wzvUU0KpggKW91b1mvtzIMCX8zk+6So6XT0KEUA+cG1PszGL7QGz2A7
rZ8lL4rL5haaXJgmRmwIj37V9lDfG78lPCM8qValPN0YmKjyKBXGckpmHR5Y0aXO
TxKM9evYC1buYdYTwNXGzL1HEZW4GRyxZd9auKimVQyuiPF7FFeBgB0UCwYjAv6d
OqzTLygysmp1QCVYuVJamoKjuP9KqCPW8lPfNePbw2DibGYpMdAU2PDut8bGClFf
ym9+MlKGeCcjh7J91zLa2BP3AlhJFrjazghGiGMTvbK6b/GbhV0BqsAoQo2l67Pc
LH8QCwetr12csBq3a0fkGFigA1+sntGu0CABmpw1AThhZufg9St658A3vu4JKIXT
WiYnoAPhuRo1Ahf7vj7waw2zGvhWpwrJ/UGdJg8lQd1GE7GWtAtZy3nI2RKwgibZ
5Vr8W0HIiF15G63BO150hcWeHQVxLPJHnxXJ/aH4UUVreTXbyJpCZYD2rMhoul0S
25ASgOzBO+YXIqbOR/AWBQBgJVYylQcg7g6le0N21q2ICqgjdX2QRiTJNwGkIR86
QM2YnECfRg/Urzs690AtXfSWQy8wNYO5Ydkl/sUzo9wlTf9vm8ABk04gtj550PTv
HGOUsZrtP/sDufW7S1LI2vZF+zIgExSXNb58Hqk3xoFLCgzYXJeSR2EmBAGNgkaz
ed6o5xIPEx8693kBxATjlskgatl64fRQpW5GnJAFokPZvHOG6yDLizRIGx3A/5l6
mvOeJqI+g1f84ZQJsE2tkEtZ2LWqgBkuFk2W8NjSjNKpXseBoaWzaaFhpCeYCaYQ
CK1iQp3ZThCQRsxmEQ3XYmewSzTl4wF7kKjw6ryh//li0ZfcbBI5DS3FIp92sZMI
FvTG5wpXyIXXdlz18wNS5IcXLjMWhd8zNpfk2kK1bh8ZgD9/HFpRxuhRQrTV+/M4
PJUcuPN30TtUnQBKtPFDuJG8yx6BuXbRYbAKo8ZFCQBkkfFDbCy8i9abc4q049k3
itmfF42jvtFH4QLwTwvijU+hY76kpLTgjfPRvVz2EkSpFx3agUCPo0i7R4rO5hTG
hGO0IsBYdjDcv6xknMSIp/vPHmCq2rLa1CAfmp5n2dHQsXm0jIzfZ2tYjKR2JYx4
3LRagBPcKC1Eugf1UKnObPBIUEHZEN7wA7WaZM0HpQO9awHNcZa2++e7loqPD9Lk
lvrq0s/4DmRNiYfy0maBtaFy5xBhzHulcjySbuseBsxNrf8hhBxKVMGRYqdatzWa
iDz+bY/jKWGSI7DUQj1JtzrJQRw2GP+YK1nrGOqC1vW2Sda7VbFVly02w0jZOMNL
eD0FJx49oKx78PLZXK9yScz1rV8YpnWV3a3Om3P+dgOD9j0BDE7JINHxeA1KXcGV
PiJEkZ2kockdlHg3O8jNFbDR/mb0A6L8GKqr2grT69Hb+jW4YFUcRtbKDjUPFLRL
yLSRpweyzn/i0NWQp0xCHbiDKgES1On54xWes25GIFJAnFafBXnegxgBfTyR0lDP
34erauP6loZzr9v1PKCwasI4uRvfPnwXEzq6FeFYw1KagpRpLaQHOJCGSxQpJKr/
du9iRKTYwmPiXvJVhp80GoE7IpvoZIgjGdPxJ8aNlKgcAjBsBLNy/20hZmYJ+cw1
mkxGEgUYPkSs4D5pFx+fGJENlLrXb6zevQMNpDMyDZv67pRiBsWkaSWeknqJ5pN/
PpxnmrE4sfP8u4eK7xEMdlxtsDnnkoSIOTIBJfL6hK5HJW4y8lIqMv3mKV8S/ay8
w+x6wK82eyoV9HvmEWE1hMkwIX76zb46t3AgQpM06/nMxxjYSUzNVGE8Xab2/zSM
`pragma protect end_protected
