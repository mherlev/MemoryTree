// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:52 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
m2EAOFynNSPt02fgV35drmVqJD/MrKXWtydJEraWAkDbZhK5y9Jbmna09hWfWSOi
DVPRmyUfPzuFk+s2+1k1Ph49toQjJZoGqmgqjFEtRnBrrqIzQdke+TN2EWJ7y14M
lyIMkh82OcqEu1S1pdkYG182J8CywLcV5vgeZ0FFJuE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6720)
DKGhsMaermxfFBC/TMpe4RP7Tb8wyW6eN9GxExzJLBSPw86Nz/lK5QuCqUUlT5s+
8JTjtLZGcIaA8DP520zC15bH6ogul5XlqUiaw/H3V1ZbgXg9TsRMI65jIJmdFR/4
HWB/VATJASiCt+NG1N1NCEBAQIMQJa/kM46lqRDHpwA5v7tUHBdpMifL9BsE4fUE
iNwIjjzsO9MvcM9hY/a+k5+Oqb4mu+awFq5LPIZpwyicmUf3yolGne827TCPFT6v
eEKKqzq9NeaThBAFs3g4OmW+DuUnM38RFCWITHbPZ0edTWsuIoX11StuB+QrPZvb
uankAkmKJyqyQmyVpa70Lqyh45zYOGVl1dfIvTjCUbc5OwLY3xuSYhkrB/CeIQ7o
hyaQFtnWo48EMJjblSLUugMJLhG2LQKB5/lsHDwamFOyrqdgVjFtr9CLTKDdNXRG
L5BzkDwHJikkoPI61lKhHCePCrbEiITgEwZ8ywBzLM3XXRONk7T6TrAIqSMqBIr7
njG3xkf7i8xOzctonJmotFD4ICOciIlDJ15REdKXQAji6Hzt0dRH2pdkjrJtzPru
JGHITlbBtFIJ1duqO3iabGBM3vYVR7FhjrdUNoswwJaGRswYm008comJJkS4HQsQ
JrZ+u9pqKAR0QT8gOONe0C8jTc2WmcSHWR5ODFFCnRlkNGDc0IhPCGakwLFT9AiH
jFgbg+/KKpErPJv9um/XH3bf/q6P5zcItPoDbvJjzNCJVymd1op0AWHLuO349jx5
I6JEQxTzqZyBfC6Hfr35r81wVVab7ClH1Kjp7WuxMWcAtqmX9rctqEr+mLP1rAQI
LsnGEPIw/yvHGy8ySP+wqc1OePHkCFL+RzUiWmGkfN2hUIwRpwni13X0sOtUET2c
szyKixCkhdeUTIRJawAA8gvoVhMF98XlFKmPtjymky899Jr5flKeH8u0+ZfVMIXY
iw15Xyin9UpUfjxJtY8X2q+EnRuOjxcXoqC9UCbtZKgyKfUshmbDmGwYTXNbGdV0
HVsq+TEslYDCPK4uA9pYRnKGExe99e2RIQgvZipR21dhUfqg60JNQHoZcMFTHmPa
82LmdMuVggdZlYeriv7w7R2KxpWUXVT7x2u9gpMBSMYlka/T3arVwYKXnQfAEgP3
2BmTZKkh8lD6WUV67IZv9p7G9eV+LE1yKCLa0TG+qrEQdE4JCFDB+HYuRz042jOW
0hXXiiiQSgb3/QBWwlWSMDTNVWqcZ0OSxac0PmY2w8N6HtCzpCsLusYbSoVZjKV0
wSvtUAzDuQbUeW/Zj540VYkrDjX+irRaxvDbt16Ynfra86lid90ukIR0WUKiJWQw
xEzGncAbYDMDiWuq+8g2Qa94QUoz7HPtpM1b7CaqRyJfV3V4Na8JxdbqALnCutoC
SF02rblTlMGorceA4h3GK5sd8WLIfLytyS93Wrj74MvZl4IrvT5RNBCjYZ/kZ81Q
a5ekOPH9NFQu4JvvW1UlRNrwSNsCKukkWyeudyQmbv8SD/noFgEobyTTwk44md/z
vqnG1nlz2Rhik2RNleuKhJVIaJXXnWXicPOlsxtgj+ItMd1rWq68QGQMu8z+n7t7
z5LQZdwdL9syIaTZEUioBMsBS1KVo+GAWPG+D2uvZyOB5um2qHqqvQqQ9J6RCw8q
DoIBrvs4bBgsGcF6j2aQSSJcCfCjnBLYpSwGRxzrGep0VmRrez5CF628ldCdtZFZ
+RzZ34oFdZyjvmEll8w/JuDzjPGIC0GMpvaZOFcSzQhDbtF8FtBFJEdQQSaazGvB
u79NMI5PUS3mThhTXVFVrEXLkblZQhQM175ipkZsDp7MqoPZmXoeIs2mzr+qOsns
fZ54U5Q6TZEQBN6vP0loDqdv7aphoYE/uqgFTeyeNqDde6+eiUNdJzNmhTZGwSKr
szfllprXsCnCoC526kQw8sFvDepooHYBv9zOuqGEnvRmoLxu6Z4Nu4d0nCXYDj3L
olde/0zk23cIYCbgKHmTh8VFAnlPeuUwBbeOw0nkSU5gKk9sU1zFY0eZcGTy7gMt
4qnGuwQ3TdzT0htWXleTQ/7vLNBDHUn/yudXvhkTbJcIO04nTlHM7GPMmOXFz2Mm
iidiLWEvYkSTLKHhfOG+OPn2QVc/C6xx5cc1PcjLfZZZ2C+wGCp8AxeCuFeu4VU6
vvsJNTNo39JzPrXYIBQmvZ792E4dDUvwsy8qw7wqfZfwEpRRwiEMlTgEdrQYiT08
m+9N8yUOwZWM0Iq4nTzE+K86E7cNi/Fne0UNmTU/HV6yNW7emNOiz5aZLHpGggVh
HA5lFG0IjuOwMPGXpl7gl9sUu0dn03jrKQ0K9f/6YEJKeiOkqhjxNW3NvpcrDRkl
QCmW81F8Y8d4smzU0egj4KAGOWoux6CJ3jJV2gA3WOMlgFyFozCOK88qx3oYbiGj
a9J7zBg5SiBSdC//ixermWMPmgn7BEJQmstwab+eHSyAoBv27oDUEmb2W2otGBNI
6TlwXtkCquC26ypGGoxDkKPY0nMIz7SXSV2/LaiV4Vffppgj53YLE99Xg9to1M78
uRK4xZRtGgdbseShfYrVnjPwybLVdrYsBAND7G5Li8qWZlA8HjUBRmZQjEW8hesL
riZjZVNjnu6+qrAh1zohlbNDX4n6fhEZbYEU0s0Bi7iT5zsVsf887RQNaIC6VFb0
FyUMkJVvSXzbusMP5vWUqA1uNn68RBDjHhK2os7n/6iEYwLHpuRj8J3YB46D9Q47
45nrzqf8zjz+alV4iWRhCBo5hCH7Obio7a8DGTJKzgYppSjY62iZrFIL/tTHsn0Z
KgHcQ//3p9RuZoXWbRWsj8XR9ecbofP/gkl37C0VRbgGx+X3aEgj/FuPf+39oWc+
l/rHvAr+ByznJvSLHSbS+BZmPMlBGMrNmWWXSbqBWZqcLutoTiioW17gLoum20n2
nUv1hwfwdh6l1fWDzuQ2PDgEo6Tdi993w/Z3UIqCpQlWLFpYoPqORp40n8CSEcBw
Tj0NGqUJWGN6fd0bVv4Y0yb/D547DkqQeOjEHDykwGGG4VeeOnUliH0FYNwuoiG5
zkwcnpymln0ZkPxnW6LcfzXVz/fGs5llMibItocU/xzfB1YTZEY4kVlFWYoXrXfd
9Kmb662KaXuK941ZBCFit+VI0N3cDoKW93m5LLBM0GghUisvhc8STpH8HRgsb0f2
UniSlV7MWLfmv4+ob31m7uosml0OevXZ7TUktBb5apbW/UWOrOEzRAMaKvmFYZyH
fzO9JRQTkWZdv7OJSnajSKMZRixBWCdbrGMurNOQuOA+zvD3Pi29XyBBdOtvNz3c
ZhTZbrkpMsCv/UIZXKQpIgetxk85H/Cck25qxKRyycB1gn5X6A1pgGW2Kw0C8TSi
wmBmVglU1KZJqTT2v9rCSyl60ZEPGXEh7m6AxCoxz1LBIH0ACDP24lqSMS8YFq7t
N6+5diwSaRs5FzHDo2IXl9RhP1MylpeD5ZWLEQoP8sO1B0kqMIJnMJ6FWY/SeqEF
2Cfz6sLtc0a2bYLTnB8YLNRSoU+5JhhcS5J/9OkyDnyZ1JvG68pOFaKBh5WDD9Vx
Lyu7EK8LI/AGyQHwl2rbzPze6y5+BuKm4Dw2BrtMYhEbL5uZXIIh2juGNEeyxoWT
PsQmfdU4pdct5pwoooIwDivMEhqqhBh49/+kL/zWXt9ECkiujJqwj9ifb7jd897q
GveeIExNzxI8NO7Sp8kY1OJB+50x9mznMxUbgbRPRGEllsUnNpzG7zYHk5dnIklo
Vk9qL/a+WfkU297JeLz4dUnA+CCBPMR9vx6KosYcCqNM1yFitZcQmD8I2umDu7xe
S2JLfZfKNDJ62+IaN2FpOg2Tfz8YQt2O4t7dXNVhd8D+RVnD3ix8+IRMt/1zQxsC
tPwtpree8/uwIx6rpoujEWCXCJcgOjYKSV1nf+TPNIbaW0uoMbkqqHQ0oYKmC9yN
SaboECapvndNazYXmxL//24XagrCXT+r2bWDnvZrgh+ZZ2os1TcRreXGvT+ZqxEG
QyCYJVR+WTYl1mUOvm4uRnhJ3sTMVHD+32lish+FGvsZvcB26H6sP7OJY6YYh/nW
qdp0xl1ftjhwLWq6rL/c+JEcikHy9HxjTEVM5JZNtVo8lRqQPsIuJQxwD6WeV6VL
wptqZlTMAeEDtGKrbTo4mQFkIzUK1Nrs8VFhO9+F+Wrlcdrjt8ibZC1sn9A/9nKL
pwPo5rku/LyvJ1iVGAX3jcMW8M5gf/c5NJASUC8JJscIEJ69Dh33wrfK98DC4c63
CqmS9esWukCZyM19bf5rx3JO7PT+S6aBEymg+FdREwq0ywg9FyekAoKRyZlQJD+W
KkCpsHtPKJVYizr4n3yLDw444bgkY1Q8pk/TxS8SpFPFviSHFYdCKbZegeDvbCt+
CA7PvKUu9Rf1miDcwyqelTTOKNEzypGyKGSRRV6Rr5SOzkEzhDx7worZFVBt87/E
CMO7gPC/Ua4sVxyXPiDao+2XWCmXVm6cuCIioihwAL0+TE/CJjcz1mg5Bo5QA4BY
1RmCFq7DEm0UX48oPp/rTdFtjjFZC63sqFZxUFiQwkMvU/kcd3k5XNqGAZ/wfyBp
+dHg0NZO7mEeQCpd6OYj/Zo/LqfNfLUe1+GGw0FV0t2bRTojvqWRsaaU/mnqS9Dv
/CosZK0UbYT24P7+VLlaLDVMFHgxsC6Mpz2/sRfZjaVYOosoW0DsMG0/k4fSt5mW
yO+CIMtTUxdyy4GmzXX2ipPbO9NAbt/o3kgnIVlF2f3L38wsogI5ZbflrASCEfa3
5vV+NeZVlMPSFss+Aj3oLsUJ5InGcxd4IlJNZ9KPtFFdiM3irDsP13gV6tVf6iNA
XPnanp6KA8H/Q49FI8sW78gx+LvG3gYCspH17XTAvQzEyub3HSepE5PGsWw7imWC
ye/0ttd5SPlsZSucUcOIHTQx9WUjqwAGQq9XtCYEQlFz6+kLFZ5KXd6FraHfKirH
++7OMENu08JwJ4YOFwNE6BwCUZTsqArww/dvxA/iIkoApZFVLrUDIVheZgfYKHsh
LcTWea4xSyVaK8zQNGIC2hvqn00xyIUsmYUxRJiwf3njUBIj3MuBTqs5mwx/diP4
GV+Gptg2/H/taWEPDCq58CGwCKn+5XrJD9HcyTVVEAj7dZxtFu44WaYclipN/PTN
TqHelhqWMQL1jzk4syPCdauBnrH334YkxPtt4l/A41RXlft5xAs3EtMRSDF8lK9J
1V0BqDY8BOF/zVm8RqWKwBnTRrCfmXdBzSXlbdYjrf3C7dH4rnBqqB0KraVGcALW
1mmXRPpG5J3HoRUOBdn4lHNi97VK2DcMJeVDcuodzmoUQ29zAzMySVID+PDwsaYM
6efc/9LoNBlvMaUSuHpjiizErGdVqgT8E0ImLBWN3zY70x7/ZS6jxRLAVrhLrGrK
tRVxSfM3d1kgDqckKWa5tr5j5MP2IQixT3LpxAL7Ro6gEcu/ZqIERTuzh9MXahzq
9sypPgHdBdmS6Ss5z9tG0MAJFuwiHCmfbaCsSoN/ZhQCrqxdX2Q6g6NHJl5DAFP7
crZoLg0wmYnX/7Q5dYxow5J5cOp8eZwrLFmuf0jg6Dh9qXgHkPvIDzzoE1VwyEfb
vB+Gz5j8lJLRzdlxF8FLxm37kwmV/FZOY/M6KIbaz+76vYQ6gaCZhwTVwOhomBuR
oCyA4WMbaRC7D52+zq88696hqX8Khi26GbgRC8Am8EPJYamA3eO33DJNBqYxodzn
zrKWc41y6ooYZ28pBmaLU+mikl80ChYY+UrKaNNH4txAAMQW8bDNGqeN+tAVPfb+
9bdIj1OFhCh6qWAutLtNrgv2KMp+/oJWcg4zvIKVLVEU1xKPxbVROHuxdQeWlTmd
OwfmGJqkr725NPZLZYeizgaXtzHb6qobtRLsEVY/ukPbi0t3/rjCAOmnLj1qT4o+
OdfRSX9vKwWsdjyU+CJm3zV7rFGB/1ZGmbq4zHAwanWRNUAKYBiCjgfncJVxrg/g
HX/Qg/2NztzyR9Vz/S6g0eZ8aXRm7GGq94mdOsWqjN1+d4ZpSonYcvYM8YKoy2KH
/V3PxmBPpNytcWcruy1hNO4Ro2egHyoqNfXbDQMMlYE2mLnwgwAykfBqBVExvM89
W7+CDFtoqXjoUrudB/++ZrMyOfOz2dAnrLFOkl5ax8A0GGyw+QXB/z879Lg8xmh+
6XHi/du+cUkyigsqQauFEwM36RuDHV2XYCMubJ2FqNYrxL4BUi7Ff3FfkyrGj6iG
e4KSWUOHP3YQyOPSd+o/XRNUNxlyASfD5J/Qh8oMwgSTYNUGm+EmZcZKmdaD7CWy
TbRe7A5/a1Tdpe37QhUqgdfmg3Kf3ij1YjL9YW8zB//RSl25odGTGB1UCZnXvOTG
oWFisUwO8uB/piW70dgbkcpnyKTJgAUhHG4a2zaybJ4C6Hi+UvS3gqY5Wr1iNFG5
EmIKeYPGQoBQIinMTh/mXwLfV0s3PGjuhN7FZOqc7VZi+06cmVqNi2mdD3RchmAn
+NnxzP0N4EZHEp2pH6aymPT9bGkkQhT1lQvJIxVE4NJBvx75TtSVxAbxLx8poA1R
w3G0t+1vwwamkGGIJopKEj3DiA9/Qr0TBYXka+bD0JAnWcllofmNMOAOui5STgfB
kDcuV4kgA69g73Ngi9sYcRaoOFkJzDksZvSALcQVWE4vU4/pookAco5Is9mtLgR8
G9b1ps74tdyztkQqiAZIFjck5gWGvo2JGTokoNPVKAKJsGxVgRb1yuH2FoIWnf2r
PqJWBJWZBdvMNA2QpE0pV42R0A3zF7mEbnv6FwUlLHknDs4vuCjaQposmBo1b26Z
63wjQdQk3guRPLgjeB2K1QZ37zBDzTJBoR3gJKZyQfd48JAo1L8rsEHhRbjvWnYo
Etiy1OQdjMX4eVaG6cUOSJ8O4mnjMjFxKxuXP7eih2VVmFQJ9xh2fHANfN78OEzr
qAjBWjrQY+fE5J3N6FWrYtbkfS1+GXmCIE7g2F2/zxJXctrbpx/aO3rsz74a+VAQ
Azy+th3Y/xX1Q24fD2CS+f6KuQPkIfA7HgZNmFn8QKFM61PnDdDRqsjnVqKMi63K
WikQXC8/BFf+dgElkVa9segJUomCIDB8FXQqxrJ2ZGZ8cUWggIOpA2kRJzx1tepw
5tTCsoescEN57SVK4vIdHCRqDBdwM8z9omgsUrj0idOex7mCHGKwIRL1GODB5xHj
c15G5hE8Eh0uQmIXL1BU4Ma1vbxDNNyYJl0jNpZu4fxVw0dUjxpn2kB/aGvim1os
AH/oPEcw/iNqsJJCsyfxPBuj3y+u6HZZrzo9XU10ZIfz3NgUIxX/k5X+V1eMNZ/z
L1xkRD9OEzg2yNxyiGr/3JRWDZG667f2Sv90zJ1iLfuDtzEKaXQ1Ptvh3wZtkZJd
GlTpG29my9Coakqvza3MpM2CXkZt1Kh27zTL6dELw9rhhC5W7ryV8cUkECRJq8jr
ll7IcnIsS9QLqetYz+g7Mi9+oVKfebe+4x6FXX7xu06kOPP/EH4MTfx7ppwVAdw5
MmonEx0XQUxSjA7kOf8cl4ZSFScz9F0NoVG/RkNPfce4Sh5lu1fKsIek1bKrq0x5
v744UAbIxUzz4ylIsn1tHTFaswZBNLZhmpDCHb6K+vk22Id/qrbmJifSA0ffgCmc
QzPvf9xK3rALLZewdewLFjxXyRCmsfpRHikdyfvgTBdtfhbv2/Oiby4jVb2q+NrC
3h1RiftnEM1hCHmZuHRZuZAHIjOhFHJy2iN7lLNU4A3Uj2Dr8Kz40NdOCwa/DPaS
/gzSDENX7ZYV+cPgl2qJmSG6mQSAWHO7PTxqYl4s75YL/wZzxZMHtTk9a03McTjg
FF3YwoXZBKiK2DLe6C6Qe2HHKV8g5HifLPAwn+8Sj9ZG7b4OTdEKOCslBAr/0kso
tvOs5Wk/huwufiKY8RIzijK2tfpS66GT5Tg/9rM6UGbYD8uQBvBPHWN9IRPcy1q8
wdoBLcs135TnqV0OjZjcYc/lKENOSXUXNszxln5+vEtHTC6+5HeGD2rjhf20gnel
gR1jt4/R7rVOYqkZ00eeQBRzEmZbv7pll+BrNKj612qzVX6wLuWgBP7S8JgSiplW
PYDRGvxIqjE9XIU4wOCjdDgPZM5Ab1vlgGpedIyV+ev8IP5rGqW/OKKQFpZRJ9k4
qe4E+exibq+XShhzBD0Ow8TPrVnD3sNLJDwWzRdZFTzlwEPoM6vBzAG8/boBSanP
Zxyeakog/IjX4EQmKE0EN5+2dRFj1iyPGbFiQOGuYFaB67kPTBsTlrlid1hC7fPa
qU+WEHeIVnWSyjeQrRrjqHtmtY6p5DBM480gCxYye0YeHwH6uVOc58FvHyAOmzr0
PyMqVWi5i1aq5PGORfsSBcVM+qPCe0e+bpNdi0Ar0LeiHv9WCUuo6iBksjrkDvDO
LZjNOrjgkE/WXKaL0iJS6R2hTEPlu7e1lxhzxetgDNTuzivjuX7DHI1tXXwnO+D+
Rw05whA4lLQYUZBzc9PWfBx98aHHWT7yMODA5WyuJK1QAYH8GQZfxeWWFyvWZi8L
ISTZtg+UB3VRpf2O4hsVQZ8+K7gTjK1f868wEpGs9hcvoTOHFMsyTOV/zWAL/q3e
JDSIljN4u82F1hN5MFqgQaSsM0HySK5a1I1OL5wQnIiaiuax/DHE4wofiwiP1q1R
UaEa8qlA2/fztG70R0CVg6X+gYgd03wL9vbOiQbEv9I9bxQqxDM0aS0CMd/YUubT
nqTe4GBef04BV8yKKBFz0oupofBL1c/bS7dj5JyoIEPIcrsWCZax0Hz02lhCTR0t
ED3+rpiWzywDCbu6kAx4ykxodptxzv1jEUYYMckwjCQSjezc3HATtNWoRWZLMLUZ
+Aq+Krzz0fvtlXQGtyuoMHb/NLGAKWTUyEM2Umb+Sx7+8W/DLCmaT1jMITTgF4WZ
`pragma protect end_protected
