// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
78agdLrmB1+YXBgn5k02GMVGxxPJI0nAg4I96a6tqLvdd6qJJzly46+rdr4PX7FO
PHDT7Tyzz5t7FYgu8h9TiLfl4LbN3Pr+3sUBTWQeQEQ85nAd/n76nNFQt2+wXy7z
b052TloKzWyIGlAhfYrWRTSNqcWHrwFEMn6uiJAWMvdbKF+8MTFOyw==
//pragma protect end_key_block
//pragma protect digest_block
qFmA8OQhnLVh3yf8SCeRTHl+oRE=
//pragma protect end_digest_block
//pragma protect data_block
cDCfi+5iUSfD3YCWvj2nczWuwly8nE5KzaT96Y/8GlKeQkw5brF1aCRHH88iWPpR
F89vclQLEXaO1fSXZW03/Ls5vOnhV6HTZVz8Q1LH5+23Dr87g1kq1AugKlAM0Cyn
Fnf3QnTpejd5zfPRdiluFgvPX4LGoVTzWnqZPPQPGNG3oOMwUu800fhn4O7T23M0
5doRAzqG4bfiuqdxMart/rkX++Z7AJNBM3UMfH2qBaOeuhio2270rnYdNsOjysQ3
g/sYIZpfcOXEeYnLtiS2uvmk6Sn1oqjDSw+iDocW8ZQ4YJZMrDq4oV24SPU/0BFj
7YGJmn0W1L+c+l5jZmF0+HxL7ecNbl2jrnKjOmDk2FHGRoneKvONX+1Ts1Uii3Jv
Kh2lAcMsp8GSCH7miFgKVIfz9P27VmEArZ4DD1p5dylNpGtctiCRfGfIGy6Nl+of
QSGmCLiTda5ftdfle9kpAINv70srmZ3LlRC4ns3N4nHpOsxsNJGXfUotT/CdOy+C
YnO6i+cyjgNWHOJCOCMSxC7MbrqfNsjZ6AG5qQztN/O2Rc6B94be8HQhqyAdJsf+
o9Mn0OrrDJ9BolUNDeBCy0RIo2ZhHaZAMsHpbk37NpEph69218PLeuT1O6cbPf7R
JJaYvuBp5e9qmbMWDRyqCwr6Xe5TOlhYwQHEDmf8CxejQcgZ80DX7hJpvTOevb9O
khr6aWQg0a0CisXr+nA4dCVjNl2VyLQGQIjj7ufCnUrsHSxu9WyAnxKzelzBuwqn
1I+bYplTv9IsI6x9q6k7WYapwz2E7+hhvrpiua4LL8NxosioqT2kjJdJ8OI1xxCS
PoUw8EKXqn2InCc1FF69CNgYHz+I5+sgBsgDpVz50ucX6AbxMYsnsGZ09/Ws5qkp
tBQvUu3lOmjPE1cX0k31PYCHehORRGN5SFMWnhTsqYgefX6eUETn8E8aF8lFQQql
hMp7p1GbNA1uGqaQ/RzGzJO4hvozDTLvxWit3kSDuJztsnyoJzgUDYLDiTqoP8s+
2Il4qe2O9S2LSpv9P8dRThDN15UX25RswcDtuEnfFFdYM4yEO6uSreD4DeiqnQT5
AHY0Q7ZuPYyRCm9dtBn1YIdk1zhZvKwK/w7HtvhPYRV8yble0xXl26yucNK8XsbF
KGyPImmJU0Or5ukaDke6q/3CGC4lxOEnYWPs1MLN+nrNtP/95iHPmCHwh1x9XvNB
e5KMrigUuLgmmipP3MoRwUH9BUJwheCXCX+yZmv+yb6bIGwu7Qbx6DN/6RV1Fh7w
yauX8aEf5fWejCtS4rcjCSmmKO3Jrz33Efr290UXN3ENaZqJ3pXWjsb0AZnfVP0g
dHRsL0i2AD22gQwpjCD2ih4X/8jBO/j5UHipiCMiaopY49JSHz2u+0PY4vbgWpbW
YWNtm5GXz1Mb85F/u+ab+J8wx9Usl9oh/pLIxwSQ6AQrbYqvDLuBF9/y2vnfHsIO
TYFdh1PKP92JE0xCgB4lU+52mk6NmfJqZIfQvzEoaAiWxL1yrD9fscVco9WdDLTH
Sz91oOwcx6jVe2WuPAPDpdP5K0pYZ15s3UHMyYJHtYQrqVm3Y3sK2NOGfsvN11NE
kbyJ41/Zt+FrFK3oPrKEBJjzNA07W+JvXV52Ur/7NMkwWJLeA0mNIWUxLjnRpthM
NVjKdK8AVFEovVU+2NhpVb9NAXJUmAGmKYAn8v1xdhiZiciuSPmrHoSNhimlGYgQ
gDxqy34oZTFaXRq3+uA7f/N5zJL/OoEllITC7lv8YZCAx4MCvB+jZKlgkNkV6H7u
IkBi47g3bdnHcBwD3KjTEez1mzVKraSYsdgnf4P24kc6wVERz58Um2tpF3+yniPE
RBwRu4M8Gupzwg51wgJRXV4MVZ8u0nJrzgAc+T7d3hxYGSHm6fIfhv9cEtlfYBdQ
48jAYlgmrkF1K5U0OBwzgxU/dsjsy1BqgRrsOnw9r7Yx0C5p+rZxtTLyW2xurIlq
dMHPGfDyuKxM72lommW7GX34JL1IT0Y0/kwGavkaRpUMh0M4ODm/9JVmiuMeIuCn
2y5fibXJYzrXEZ/L3Hs1KjVeKJT2cbGh74UNBIdEE/1D3ZbWin70a6jeacBgeIAN
FplnN4aKG5pfR1wqFpTn2VsCC2/BpgKQQEGf4yhrbgHyv8ICkhVNd8niHitgQHDe
j6o+NqAfplsw3v5scS1//qHWSePajRfe1JGiC2qOmvxlES0PJ+Nkl0i7hl375wm3
iprlcS1s63FbHILFoptZPaNziZehqvn/E5hmJl7ZObTReSfvIPHFz/MKXNDbjdBs
AHtujlaMcGPCP54CCeiIWbN5WVBDwXxqN3s1X6PAG8GzFLzfyRtM9FZfNAMOolaf
L+snxZAtVTIVYiFQwgch4ltW++oOCZXcYb2XjwRkmRAaaaOlJi0z8Nt49H8GgPcB
QBnRh+DRu/x09ejrIm2D9EmYYcQLQWz2gWYyOOF9P9zI1SFb83zzgEEo2/XpcvM3
Pbm7a7zgQ+8KCejzKH/ppct9Gh6GjBR/cycG732pWBvtb9NqtrP2UOGz0xfJl/+l
l8LZWpHfSmlXs7utoaj7bQb3CWiIqsdaq5g1DuaJNZWxNSVWB7LVH9waw9OZUq98
LJpN3mVnL/6zkAeShux4V8wJ4ALIZGUzULafGQcAaWCfPjGbRKP8VSqqELGDQq1p
w+f8ndUm+NMFAV6kYXOxTzL35NRs9nj/BLg7bRwmBd2e0bFYASvwjS7F+QLxiMBE
0Uqw4U22j7fjoCYr66T9MO6Amv/NQaronRmrGCygkC1qksLTi6KscqOT2PRNx1Oh
lvNREWmCBR19vYuzXTjIiS4f4oCXgeh1Pv6wbtP26Phx3aRCaGHigFcXn4Lu1OME
krl5GTuC2fIPu4Uwaq12zgyrez+jlZWbtMnK90NOZl4KKwRHO5L3TQJBZKKHgTQ5
M4S7EqQTREPG0lSZkqaAgsWrShFxt9X+3y2eHypmU4McdH+qQE1REFmqXmHaRfge
dWQWh1XvA1PoDPJZVL/A2IGjpm4yi+1c8+zqs5TutZ5muIfEw85jSXLD4d0duD3j
bT0AfeXlp0ZpNt5NC3wmZvovkV/EkypK78DhwGEgM32QUC1aBpg9X6qNrsk3Ft2Q
SdL1AwTiogtE3FVwaxlXIff836p9MMpxku1+GjozBg//SOjP1+Mod0zdW34u5sJu
bm43fUfg/woI+05C+gYaB/94PbwB9iFcNqvgTqlZogmqydcKSivM53jg1AfQS4xx
WgTyMATaR2hcGgneeTeLfCHInDw4Rbgpetr6hzccPM4vsAcLZlVaxg/Jnv9xUGfJ
34fepG+dVYLTOIhuOh81oaJbkwQVkk0GXNXmbX48MZl8bv5QhUkwhoE2GsiLkaIn
bqQVMXSSXg+GriCCbtC/5BuDagX1IIKkWw//K4BU0g5dANJOeQr5BnWDCAYkvr2U
LovN+5f6qxC/Cs3s4UPT9XnHprHhp/XK1CzF+Q/KugRzjIkUpx5Rf46CuBHr0e9p
yUYkJULgldSkS4v6LqGnd14s4UK0EYW/r/vnwcp5uudoL3bAY3OZ+zM3l5mjyxqm
3gbkTChzvr+rDZ/DveZr+28+K+RNCiN0zDlVbdgC64+Joo3Rx2CVS+XZnaon7IEM
UATp9tbysiuAc+9eyREaZVK4M+JI+WtW/yUuasfohERQvyZUqXnQ9PzXD3uanQSd
T4qTJU0uJMgXpZrHVjCtP0m3vV4gZCSZkspHe2mCkv9sd2lw0Nm8m5ZBHO/dM1zZ
wvBRgbKvymJfkZGCjPSzR6Jtf8qLsImlxPpxeInltCfQpMzUTTD3xUwe00vsh35N
g9PExEqvSRCuDf9Ni6/zPpsyi3Rrep/8m+zTX/a01y+ZR/Yn1vOmRHMOcHzLutsR
KfX4WIW802wu6+muR7DHkV5mfPw0ajBp2UoTg3joP+35ZnP7NiplchyiSrtex+gY
ZUhbZddrHiHbRgNbvGh21G5mhfLMtOQRnRuAJESOrpL/NISVFisaqK+klmmd9I72
5xJeI9AdpdbPv+bMhb1cXfIfYCJLadOx9XCo0LOGj00MZHfsVtIN5Zue3VbX36J6
+A+VAIrZO/5QeRiK/LUZlM0NAX5RI5aUhewX0hVLWnRCZC9Xdzlj59v0UUIva+PA
+bu9+L1EABjMsM7vXL4eN5VFouY4FqnmzkHM8XtHdbhmcYpZ+T+q9v6riKiF/25k
jn0Zoodb+1df0/Y01if2EPqlLAU7IPMKtFsBXqMtAjVDo5bYv5TO9Qw+PRLEl0Sq
0BymCqrlNiuEJcYHb/P1sQGYLOaykKFxuNFwfkQuuP/vq9xKSBAXQ5nBrLjPrtmP
Wz7836Ozf+JUiQPFvZSZI9YE70hPiOcpCVPt7SZsQXvIUfTvBWmIy56072SYhKph
XmhBp3zZk59XMrwR8VClVp2viR+yn/JAUZ9q+pxdaFiXeJLeN+R6hkZ4JDginlmV
/2TRJwhJxiWB/U+k6VyN+J+0W1uPuGa9jboyrxj3YBgnLSOGMkdnZZMlw10mDSgb
BNXWh2qIV1rUTUIwGmJ8ntYJGBDkl/gGICHSNwucRYjKP6Cj0bFB5jnNX8iJx7D0
X/RT5hz6tHfnUcE3YlrFd/Z4NyW+cRw+xh8xtuxG9AyeBfKpZr+e5d8U6EXxLgdd
ceRIvTqmhrYfROIOv56TL+flfsJ6AcGrZWTuKDyme6qOqb1Pm4donCz/pQ4Ahv2B
0cKZ+Y8BxOvsRJtwm47AJbcPNb8Fll8rtTanD/Nb84UW6l75OuuQuZEoDiTmI9ah
gycpv9vNlH6eVemhB23q1TttBXIQMFRimklgKw6ZY89XlZdX3NNM8XUyb9Hb/rqU
PEH+wxVdg8zE2DiG/gRWZnaCT+T1UxSmgSDuf/99OPZ+aMlUGeB6zVG+QGXIC6qJ
JL9/LxUOZbyunHLAUCrF8r8Ju7CtzftNrG/IMFsYTMOKHQFjmoW+LJP1oSi7lLR8
tJ5p54kkLc5G/mMZudDdg7WEGSDCma22kqQ3rz6kziFNTfN/UYnyTlqzuSZdBRYN
ZJjUCmEIRgkgLeAqA9VAqDgxlI1KVPOggkez/SXlxwEUDhA0b5FSJsdzTrftSndd
M8sKO0t524JI3OOvLGnVdet7s9I5YORZsD8nVS+pQfyUQu43HT3Cuohj1jEIMHUG
Pa9m24rIEV0PnfTIADkML3ccA3Hfyf3O6oY547JBux323+tPq9aTmoDIZo5nFp8h
ckuJLrOBxfbcJRMzYrJ8QBafDvSQbfsYLE/8NRXGdA6O6pUD+E3qEklueQOENwvP
P85Ar7ioJqDyv09HFTlaSQdl/msbpYomtlcMTXe3sMj+GVdJJhjCJLXTdJjY5z09
K71Sr1b27/EcFFYZFPlX2LRW3RxMT4LtyRcDHbajt4OVpb2kt/VjbQC89YZnuuTg
DG1M9kRRsNDnHWLgUdcyVdadZ+Xj5oz/1oOhSvXwyspePDXkn3sCpXVtJreVknHA
BgFi4EU5IRAt2jCnxVXm6q2VaN7ZQzHwkHqFgMcsBha8XKjj6fvBA/o2xOKpiXKP
sDEbEcpB53EISbzJ97QnsBMfDB0ZTBeAMOe/ud5Zp5X6pNDl22vTxlDBmulRDGtM
+wY3l4PDIhMXmYFyfNRWmBhB7uMKEbnIYsjdv9ghvv1pb0N5fZJrqi9r2F8CUvgg
5mSY54PeX59aNY5F5ZBcguR6E8iohi2Qh8rbQGu0wOchD7OyPB4rRUQsyV0BxQrz
5UzUc47LpHPg4hhTrv78/KyWggzmUkPODmLxu3ddRep74FzTi/C54aALnLG7cE8P
nKxB9CrIeA3Ug9OhjL0SKDCLF5+S/ZAwb5fTQPC2rTkhLzxrxUcqMK4GAl9DTLTM
yNazUp2TfrUYttrxuPOYtBBWacHk+PUqzfnrazXnnS+5hWvG1ZZpG7ujoskOiG5y
x+kW6nu5nHPzFk9f7xAUR3lDMun/rfEdGz0anf9Hj+jJtTt+6vu9nsOrE8tQpLyH
Vfgt8A6C3SCDzyjGHYE30hVz89yRb8dV8yM5d9Yc2sLQF4aFou5JqAU+/l86ypNU
DTr93XO9A1dBrpvqaQP9Vj2Szj/1qF4faVPS4forIZU5yYA2V4RGZ0zf6ojM/LGx
CQBVDDdXrQu+4vrXcrtYkWBLOOC+PDXuJEm+qNUBUNecm+k9Vz7nSKWg9N3jfwJg
wgkhfwTB4rYUC3pMNrmwSp/yTlcMVQEQUCtCuHnc4qyNUfKtQBgSWnMKr9do4qB9
9WZFORl8PlmHodvRzoU0BiWIQ7HYsc9DaOiLgqThD04rM9JR7IEoMu6fu5bOfPMp
Xx+qJCw/zIV/8dK5UHzbn82UUslK2kh/vY6Y9P1O2GkmmdASOB7umK+IoeqbJCZ1
Mq5fvOTZXmRFblxuYEb2wWBLEyBeHbLawmjP+jrtoHxXZJR/b/KoABQ0rZExQdb8
HUT44aUqgj7OTWL2s1UtCDyCOm/weYpiyEVecrlI9E0G7zPYcZ/ttjRZa5zSsDhq
p0sJ3nTl9dJd7poQouZqRvzkVLFSl8P24pUOsfNuN5rTDXslDysYu7+NaYd/xh+0
lOMZGBYr+gn8p8PY0x3bTcfabAhuDpiVHm9VrxY/QFLVZiUZWJzbqCeHltj0Wcdb
Apc80a19aAp7NdlzehcWwNzwNRyF+8zHPbeMWcNQmQHMIlla7U+nxTy/dxo8uQ9o
YkscY0aKQVdkGZLkNk7awf+2uxo/EhYl4/ZPH+e+MMwCx40ZnD8SfHpbo3xJunuM
qNQawrnldYoguxt8Es9Fn/JkaVwTaHW3B6TFOD7joT8Tg1/kFxR0coJQD0kOGAws
2RQcDFtTm3T2CBbyfB9ZhGJGCj2cnTaEa+nipC/kIzTxP4u/7ctK2Fi01g8hLaUp
2Pbf2f7apcaG4zszquXtWqVb7+CSwHM30/fMYS7NjoYRvFuU7C0feyXdY7S8tPc8
K5ztVdH3DOIwbA+/m0bMrohCpGpzxIZt7wWz16XqYCP/7gOFVgW9lEoMeMJn0Gpg
le+tH+lGDrePy4ZNrRk29SEhsl4fhLrhFK6eicbY0wJk1oxhebqIqyawWbNXM9Ds
UKp2HeNuriD88EGLqhGju7PQeF+zakmeInzpXZHS58QKrqRqDUmVgWGxcrq/zlZX
i85xWEbypk+57oCjA1SVshVTz9RoMUkwNLfztaCcBAiKlEuRd6jZS6//2OIZ5FCA
ErW0P1z9kM20cuOwjsHB0LKME5WFUT2TcS9WdrvLvOZhGaPDosYUEY6uy2BUbIN4
FNW47PEooEsndMZl69lL1j3isM6fLDyqT0PrSlU6jSqX/nngJwAWSZzIoRm62Hd+
GKq1iIr/MYuuJfnry5Wvw4rM28h7rbAYM1nOSr/3oHR7yNlafBDfTnGfQRSfKjAE
RsZBRQ7yDfbXrUmmuAUGttxFTTKNO+YNdB35RsJnmKzPz+1TaaE3RredJwmT/meF
+aVe2jBk0jqGMMdaF5EurEsQu4tLQYu8hwH5JimAqb080F7g958dDs/X8BrQSysE
PeEpGe3oD7ki3PzqYhSK3gyoAXKTita+OfXK25jFawjbxjb2ktoxjBQkpMWmO0Lw
jW3rBHtlQWkRmYlBFXRjboqfz93yFcM8MBys7l0cHpensS4cuiV8zaDEzbIhvqSg
9Hrc+Bbzw0LnO12NtXZJxZTxa2dPUaZsQ7pA6ot8W1PTQi6PK7WlHf8bjXkQQOaj
xOpy04xC5AdhkuMt7BsUxNn9Om4QUTQ28WSToKGPlDQtIK+BBODi36sIw9PiufNF
S9fRzDhOEBnzdHDVdX6v63BYPwdaQ4BD5/FDeTy2Dasa3S4rnb5O8vikaduUSf3s
Cgsj9+TRD7V5Y+rSg0mqizr3IP0CDRK630OBNpWHuirvGdGzBkSm9rzBbEx7IL4p
BV/2H/9mJiscTei11N6HnEyvohb631hq1n0MqeXhD3FNBEtULj0JnFhatCz8dNPs
PXjUdhwQMq8F3dM6+XlkgSXRKlZ+bDPe7rvf+J12PAV4gyCu31jE3MjbQ1XTJ3pK
2kYqoGemCvh0lLdbVDniESuFEOK71aPkD5mPssFf2KClwHdhCZWW9dVuMhL+PP7E
nZIisyP4CyuodwFs5bbqgcfTmsROA210bUZHYwg0QfGoJee7P8NvrzRcKFm/fV7F
qFxua/Tj7t5MtuMFVq/Xmr+GAOvJozCyW16bp4q/UcdKY4RU4uATMnmtylccREgI
wBpsnT7bcjkEd4Xby6WGuDh7kyGLGmSsDTic+K89RUbZv656UhUQ1YaRN9gZYBQm
CwDDwY8twDoXsTtCqLZHEcfzD+DmBkOqGMj/VMPMpkKNyeaTSrCHBCtbUtMUtmSz
EKi2kkYhgv1K5QkXePG77EnP0Lm7kLqHIfTGZSmjqU4son7kNO5uaEg5JNB7X3Ac
X/H5cu9dtJztb7w9HO3W8zkSa2saKlYKAY4wTk2SCk6GiSgrBUFsJSl8JAvoUFfP
oOk9H/KC0lwS0ifa44yQJ9movhhLZF8pVyksjVrr98sNEra3fRk078mROGHjhmWJ
w3yC66TUs9SvKepc2t2KeEfBguUp+fonuRsBlve1w0/NAQB+suKGJVySBvnxyuRm
mPQW7p3cup3OdkLmA4AvPAQ2AcmlWRI2Jjc3PqzcnDJwkhbvLAqSNDQxdiLyrGJY
/umn8kPHOfgBkhcoTPHNf+buyoCsz9dPKHHwxyVhEBW6GFfqDd8JKhdKKBsP7QaC
TIQhEkvKHyn1zDwdMY8Pognc9wCadPWOHctM9NHxq5cJVkCP/0Ge0bDhSWW1JfIw
RqVvocaDolzbe5aAoG/Qs/Daz9TOPeY3yE1U2NrRY763OKj4/YA5Bb03imMyC5lE
FIWr7Judndd5hMGzWMXKWpU4ix8kSKzMRdlReD6zxOp+PS03VnzPo0Kn6neINuPb
jE8hXQqypSHFM0CP6lVqDvWw4DH1OEGZbg90/UdII+/Aps+IgXVRMVgNSRjb5VTM
sTRhCXTyaSOgMWxWt5la19RvISveUg29EylpAK7A7BiubQywEU5NJ+f6eIV8IdXj
+Ak1rlxmAU39mobPMy3APPh6eSGT3HWMAINy0gCcpUuTmRIVjsHcdS1JownBATcU
KRXOioTlwW32MV7Bvuq2/5sQkg3ZdoPFrM9JF9R1hgiKxGg+j0PFR8IZMd81winM
Rx0gy/DlTHikw2q/A8lJ/ericaERuZRdxlZcTojeZl8tc/Vr2NGMhM4GR826cCd+
qz7X4bJxSrt6ZIGHd7SQV1F7g6EyCkWKV1YjnjXwwKnvMODk6YB+P2FtW/NRp1dM
0gkS1I/yq+0pfRBZsUOM4GBRXXVsmbHJ5zhTqVn5CkBFKDwrhI5xJcOKJaQw/IxB
PcC9ZLEQS4prL6mugnqJiWw9RRdsbRN+OhT78EkICnEB/A8IzE9v2V5+k5F4rLCw
i4TRGgG304HfkrrWNucTwh656z0sVRzfjGFi3OSknAqxbHe6JFOI+pMBQ2uFcn9w
XHWFwWHhrbuOQD2EtyFEd/1aEopSgOQ6nYF3diYVs8WPc4A2F5jZDCfKSHpCFEkb
u6VCZy7Ym2e15M0FaGYu3tnWZ8Y6Er3PEG8idTRz5J+RHIlWrpHnCUnvH9+aLjcO
sD/37E2uQhWjvegSgh9xOn5etSeAiomevA1e1ybxN/FmIOKSEhJkzkguMlDgh/z3
kW0DBXTiHZW1h7pfO3YRz6i8Ug+whwEWaDMCUwrMS5EWn7EN7TRNxzwE7CvBhXBa
6ZEaGlqg4dv3XY6Sp0uw0a603q0xe2U9pRDW10mfnOLYjTgTJuE5RLZZr54Qbcda
NWWhrIdgsEkDCgDJWbRI1UIemPvgRF87MT8wfSi2jSNhIRtu9j4hw9EKDpSH3oXM
qFkjcH3W7urTMrDnqIcGmWjuuCdfvupKKTYslsED770xkzM/aX3vqPzUSZBnu2D7
pvS8MqG1scPag1xdrSC7K+hSnAweA7TuD+o21U2aSBRjzywpfYEOc0TV9OCvTYaV
yyd/vJLEMzkGtDF+EqoFoZ6dCvdlGqxqA/jUVm3pUMi6UFKTHKYBQo4ZQ06LzOSE
hjntJ97WFfrIT0uLAZ1U3ei72EG2XPm7na7FBIYmGDanf0ENPSiQfFn2aHxI4dNf
0ajGLCy/3SQriZy8bVKXyZU23vHKqDoXxN8SV+g6VWecSt39UVoPx2v6nbtzthuL
l9FH92NKM0IWu2GsWy8CsrzZ48UwsHz56PFCxeAVjV3PNk8f6QqVt2EGVSsegOTS
otY6LktPO/fCigq6f+s2ZRZI3zARUBNqF/xUDGy/jzeZ1F1oztrlIBtrrv/JGOF9
mrOKFs929QhTXW0QJMBezZjnmnPWdoVzOky4TPNsWtdbZhG6pxQ/FlSjxn5+nKqE
lFcObo4msmnJ7tZ+uWGT1n/kME57XOAxdiqLufxIDxtHZ5ouN0eSTl6OVppjWWsR
obV/0qxcQ00Id16qqbchlKqVZDw2padMmzeXYQUV/kCOU9n1WkjyUTE8CyCuHD8O
ef52vdXy3f6UOtQKQ/zpgvxa1FqVaglcjcwU5fYB/Kw38vmKKRXx2G5TBtUnVq9o
Wn2PfuargMbrfPMPCmpkADk/Bbo55ph1r05vR3CzQJmTfFn2IVnuEXAqLNYrpQ3C
BViZN5Ue7/9w76RD9h2mdQbW9YNohs5Eh/s4YoG7B+XBPkg+DIlaLPhM9WeRSoSL
fUCyMvb9RQIriNc9RX4PqIJ6SERMH7Dr/JexMnyooWzQV3nNVE/HYnxIpCRw1kjI
OldEVzKKSE+zAZqHUrqFcaOZMh/4o7cGaOto35fghx4gaEdKdVOqNM3Ec6EhKyP4
crNPYzgJ41gssgpOUmgzWzMz/NyGb9XM7uUnWhxShkOR0+3cB05Q5WDDApduG+Og
MQqTWrENuTPdr4QF/rXpwPgGL7MFUHniOvPdQR4OjITSDtuAjdoKxZRtwY0pxUOh
rEi7c3XXtwf6XHk3gmax51F0dGaPnu7d915BRChXnaut8TIFCYUeeqLn5WFSu7y1
vJFLCDpFFfh/7tITUQG6J4RSG7BJr60HNWSMIvg9ycJqaS64BdU7M1AgZ2lEjYXI
tA31AAfPo07PGR+nviou9/G+C1k8gwGe/xpu8+a2ju21LFDvE6plcBLb2rE3pMgK
bEwkOIF/mdNjhyPwg/n3ZYbnk3HZYkyD44XztH9hrmW5sxKPlRvmFvnkwWUqr3gb
5Ex8CrJIl25W/2zp9Y7a4Q2Nm10JZsuPCnzq47vIjdZlVTZ790gOtBh4RR84Gohh
K3FXZemoeWdLl0FBrhdmkGI7yIHcy3tjbV5Bp+58RR1ZD0pi7iedkgVJEMpwNB3a
qpTitN4IeT9S+9cUiBYb08NEQXVtRibX7G++jTjfq23XCYVSHANdnrToSxcMOYUt
M+nB2DbxCIusUoFHK0cHdTTVt9uoEc8JlS72A/wBSr0O0fA/SAxzRThkA8YiuFfX
7rpp/CQGRxqSooJaQrrpX+VbqJh9Myd0wQ1yyFx7FtkSBiTAME7u5FaSZmI7XcTe
1GYqQeRBuZzf6ascYkZtIGROma8PZKQv0vVLLHIy86DnIqrVpuVereLOAhyegw9C
o7JLcDiZIT7I0jZs2cdbmMQ+gfwxctmouL8sxIL+HG8RDroqG5VuA3ltlVn4RGPe
xBY8iDgch3TAV+CH4NNqcG93rRIwNICOTRfK2oFNkgM8/BSNCUlpob4fy3ASweNq
UIa1nsQnukuqYK2tMqyJdiHc57gYQyE0WAW339cvxTQmIYbk1lHhUQ85zAt96+AV
tN/kkqBQ7nR3z3BaZS7D/qUBrmtcJgRdFjUbW47T0qeL3cofPpCOr6vCZsWO/rXG
+ftLy5H8NysTpE/jomVzN+NqAM4JrZtbe+ExnS+z/cozVYyQi+8V+pnHcAEnNTUI
uWWJMcRx0XjgN4E+JsNTLSRN0Mbv/lFRu8qJ5hcJVJETBpnSKvzhSjj9zPAcpcfm
yWHMo0duOuBPKqMvNdntgtJI5NLgDuQ+mCOP4KQDNhRhOs0MldTAcTk6m07UBEed
t6M8I1d6QTEOUT0BTPGzlu8y0Ihu3Gg+idFM11rOFP5Ccdo4JHH2YXSD8SKz1VSD
sjlsd+B2G2vAOkJoIyg504PJFT/kXy52E/hGgYv5TCIsFO213BNq5OHZuoNxc99h
yPDxOql1+iOK4SNsJG/85qHZM/vewGg5l/AB4q3as/Zb/o3Z9BB2v3M3tovm0719
X98DfXcLeVKjX7+d1j/NMvEvHmMHc15sNPyoB+r60Ak9w7Xn+1fAjFtAUi0bueMO
Gs3hPQtaw6QPQMvGvi8c37qLaunEgMCDNjbxqsca9rN/PHemsime1P3V56GKkd27
+EjuyCx2kUtYpgk733MZ8vXASyWlJCMWXydQ9zSRbfOp7xLkjYRahk/Aks7EnGc3
OHPK6GeR22jOcFmKmygbg8ddV0CDaM0x8ttGhQHt9ooVjU4hSUcV0pX/njySr2N5
aKobecnOqxQFYCFKl1HiwxjM5zjT/nG7q5IAhM2jekA19UXDhAuOsgBF9zV6PIei
vw1baZcHwF4cmJKfBVfeEF4FKRwkp/zo3qRn8ws3HwMmlzXXcrXGEccaTiJoh2cB
RSzgb46LUjDCaqyQ69//4nlEkePBnqRGtBJOG1QaiYeFlt13qypLQzMBGs6IjZqH
RSHQiJT53JhWKX5PyxGgOYUtqkr4mo5DtEEjca0qUK0coz5nYwmqcJFtvgPHTnzI
CLz7XUmST0In/8CRNvTtRL+o8fxSgB5sxSEjeKjCn1uQ/Z59zu/Upic7jGeVxClL
6zqq4U/8rDZGhhCx3XzmO8I51mqXCf3ODttDkmZUuGB8k2BD2beHDmxVyfLREac4
a3DmL1cZOfIctGCeuhssqf7WsufKfZxioKaa3HX8AIW4kMSlYk+OpG1Ic8wwaWBR
k1fy8+sjlXtvNQo2lQ3u4pYzLBhoEvrDORSBsyt7YtYyeS1cQ+stKx0PEJaTalN5
D02i8pSlnI3rINmPmRuVnJjvCXP1RscLgRjTg7F2/UUqLQnuDCCpOT5NK7QkwmfY
3TiyhsbNv3oWHU5yPfOi3iOuwpzKPdY+jiDF0aemi8VP6sX92/MpBA5LucaUNXGA
bo6KekK5Hzz8inOjz9daOmfVCVseGyl1HSiR6zUFNKRnQtLCGu1k+FLMrtVC00xv
FXZPTrEfr6YB6a9VGJ34ANu4m61ZxTdG8HgfeHvQKiIYOja17kS0+2WxYJy6Y9m7
Q625MjbSQjhX+NDkC1KIfxMN12hgvwE3NiTsWBZaqLHWXIx3YVESi43ZRHJzwFXd
BBqitLKDgDAA+5W+cubN1OesAaw4y/gYyiecSOSj1qvI9nOL/H86Scg9GNR61aPJ
2J6leZ7pNKr7ekgSvhE86gLeeL9Ol9M9PelqyiUxHZWje2Mj/Utw9qnPn3zWOEdZ
OJyLSNHhxkGEYYTBDOlSV4ux+jKaPxLYj+B9oEFVhr7xqmTmHlX/IwggYI4YswCq
Nmz9rJe9mOPGHi3QBdX+dxBMliDUt3bPUCJ+cYO05GtJxj2L1HtO754OzrJzs8W8
Ja/GXiJCtAbqcFhqELnYjSiPmHxXttb1t9I4Ox730dfDvOA4dsIKdQdedQ8xz5or
dmTeDsXTaAz8K2geYgO9QOrVCDFDsn9zwomZWZdecJA0k7Cwg9aauiLYlzXuZa67
5tL17ptjmV5B9PD2SMN5hNcbpK2wa87hl2ZM/1DiF8CLe4ZP00ROxJEUE1LCA18J
531ZoNBxjWa/Iabw/wazMDVfc/bOxmP6vbs0TnHZ2ClhxiRqw74CEjgX02D0/UCo
2yzdaR/5cVOwpaRu1pA/ZoItubWUzPE4llfuFyNF+HPP4G8TWQYDHAdSg5kjcFCf
Aa+flmT489ifXAHHzWfPQti7xjkPtfUz0G2kiO1FYLKoHvthnziawQmcOPg2GQJ+
fJEU8cwVTVI6zuIqoYu+tT/4PKudCUQ3mbxvcxk6R4DnrWTke7BtLAtNYqqWj8Kw
k09YO2RClcb77g7zDDApwen3GcXd6VL4JywGe04I/f4XTfZBx9Ln8V8lqcAmJUWG
iN0wuZiLx/MVUcc693DQncUZbqf+t+L7wTO4veWaZqZ2cgQUaMy2TfVb2xY/MLWn
MXm3xCe3miXgwyPanvxMwhVbcbrv8JxpnaLAytyyAqrvf/cchsCjwj8Ws9ZIbJHw
3tzxWn9HF3ricioDnQvqmGeLwpuzOJkruu7z1y/AL5JWKq2bSIJnPXrWZXwRl1QW
3iJjHSFfy/HCRUVR91K5vyNEfy9qDWPGVRJHCtz2FH6dc4Gqia1O9owPiQYcCe/E
EiA82Zinl+L79LIHo9GC4v9xwMUJvscNcJISqK0BJziQWhIoQImY+Ltmsd7nSCbK
cbUwSbQOKBOMrMFczptV0wWr/ybEe87JEsOKFl7oCEjfS4mO59aTS6cPRS+bQnoA
huclu/2iQa8tGEl6ZmS0szfkq2GeFXyEaMr7oFHxK2VCLgK1CV8nh9f2URcOAliR
dPP9/4GOoh9CE8wayW40ZuxSSVBZTzzXfBYLQE+9xz5tOjSDOAS6rrfvzNHkn5is
/H1CpT1RU857GxJYTLe8rsJnT+4t07Sgv5h8bFSSnWj3w0uId/Z+oMjRjrGyiYL6
CDNAuq+tvacKilkyD7jtkX0jdksoVp8MycBh+FvYOzPg3NmnIhM29LldJhRLb1mb
8YL2B60hVZa8gWibkTrAytAOoDgW2nfbkQBqfDRLAzxiwhEX/JtAyuRurBCFAUYx
bZDkawURQTCRoeJbqCS6VRG9bLgn/4srxiSEmb69xb4nvaLFdNVADwycaNBN230C
1nYToefvQcRVDcCmXyWLfpauFYfb3384bmp9j/+ej++gtXyJaTvUOCs0WwkJn66r
FOK9zFHzjuN8vxXgFA3xNqu/DvR2vrLS5pEbEAz0REu7UJLfs6Y/8Nr52gbomrDl
8bxK+cRJIYxDW/FOY1/54BKe7eXy+OITkvcPw87Q419xf1qC4912OcPYygudiFMB
1giLf4gJRzOgbtysrO6+IAP61iX5DR+qyRe8qjFcCt7geQMHHmdt6bFpUrCA8E/z
f9U3IlvuP4TuoJoivDo2A4vqIO3LZ1LEJi0UHNZ3IkkL4mVlSvB4PEGVc8t+QR/a
JVXnqxPSnntjtS+vhFolTFI/sIDkVMqma1lzNNPVST8gdFyv3FQD7cqXIvjrVlOX
+joZOM9IPQa2ae59Cmf4sTPRjPswYq4nEtiUGWqr3ph0JS/eT0OobHFt4AKb2ec2
k/GuMhBUWCDPAsydPBYKilKMMpxk+zjQxOAExoYdDZJbERcT4xSe9Ie3ac0+dvDk
NZHbpzLzzbYMgl2HVzTDjKYi4X062iMVCpBwxgyEzsk7QIWiibBS/B2+fZ+bmNU5
IxVB9iwCPwq8g5ioFMR6jQJ33o4FXuJPn/mL1K4gpGNdBegO4Br50RXqNfxOI+ye
YPTd8UyFrrAYHHLFCjW/J2cCM+xTppIYH4K1T4Tg1ZKJ4Tr/Clz4SVq/DcwKIFFj
gKINegROgn2WjoTrvM+11/FQm/1EUPddijmyqmPaaxnHmw2dChgGER4l1CgOZ+2i
KnwkXkz441tqIAw97fK0Hn0/tdXaYPAPa7M0WnlOAcId5Fm6PFfNcdaTyX3pktIR
dKl4RAOkLh1dwm2wCjWdq7R9leVAFe6tNIvaMIMnRm35AfhANAsl5ddcmKqfptaJ
6cwJc/oExU7orEqSvWpoYPxG/zJQ6advJLLwkDjaw/PGKHLxDXn3glxI4lrZrKMG
hk/o47A7actDtBo7Sc2E7eGBs5F0HmMGY/5n//jk/XSd2ZWUSk1CHuXzs7QN0Oye
fN2V7l+MaSRVBufJhCM+W4CKjpXyvkFDlFx9RxC2xoUPhs+W6caMWWdkOh5gJ67a
qoDE0B2OvhJ3Gtntq9iLkVhGfg9LRITlEVGLFGMD/IIonN3AcVseob62cswc2e2S
HsImmXrV4aa1TYWsk31htYwIJ4jiLXADcZ0aY62+T5NUplibxq766Z2pEey+1bPb
RTUtFK2ikpU5onrbGitXvsm4qUJwKZDBeuRwjx+AEA/7gkvCTkwHSKKZjVtOcLYh
hv2v/22CIoEtFQoxxqio1VETJ2GUz/TtpyrGwujQLl7Y238tzZrxqYdW5Bo1oVxn
jiXtbBW9O0246/jTpzHt6c389BCtQfeztbSln50uSi7b/adoCCnsyrr/p+albueD
4o5cUpmHIzg6VLg4xDW6NPkMt6wkz+QaPkJZKly9lD7F82wMGsDYcKmK/FcfenDY
eztq/NjPVSO1BdFsEkhCzqcdMqUrr/yNaQ/t/DV0Ui7F+qv3EmZ73FTvrptbJYhu
YwL+MJgzPo8OkIyAApMAYiMmXylkGInFieKFVcSEZUmlif2VFxf5TiPebZ5lJdiD
vRnInyHast9gpCVx6gxcqwE+UtRCQZNb2krfysdRl5iZiusOVZCMuLbF81TD3Oij
f5IP95+JCWX7f5jahPrJbKzVzar2SasxDLiTPy5/Y7zML8pYoH/ynkDNDfpPiJgV
KKMMZT+O9cFp7t+lOWFulrPBVGxlhYuAiku40urzrqyHA6uwxKIYXMGPNCpu8xp0
ytMFhC+uj4BELqAsupx0tEVWvoGdwwvoBJlwdBoPeQKrh/kRG3tA+Y53Q3KDJ0iu
i6LI1Sx8J+F1bBYl2mNtUix4bPfVFlHm2U6Oe61QGn4G+ah54m5aIwTDP6pIRDEV
4+5Z343WKUbhlZR+Q7euX+OFAnQQcp2eDDmg5z8BpYJV703u1XhKs4pkhgexuGnA
V9pEls1EKyIYVRo9bmlatYes+6kI5cI7c5pnlnXtg4koLi/5tFwrg9FwaIL8Mj/3
VZZwbsE+ZcoXGWVQN6lW65lnr29/pXFrCimDfjSLsyjEwOxGlWBYrP0obm/yrHEs
WlEOB3M3SLQi0NZK4nTrafDPMzTw6uosntUMCQC5SxRZHzBXwJiooXe7ClES19Fm
Obtzw9sjka2ImvMc8mGlJN0VOLUp4WXFuRmv+YjdkB2xLiUK62rE+NTJKAn+q+Hb
FMII2IfW6/z4gTWp9vqCU6o7wSaOXvYHAqPaAxNIoQrnWzFSWw7K1Z8tgNYEmAPm
5c36zc8xl7kvTrLDavRKXZiYcN9vEEwtHiU/tF95+C9yqWWRuT9RHT+LqvGUGTv5
nZ7am4HtU0mE6tNFchH/QUHpk4vZ05d6192RHt7Rx3B9XgdxwNFGx5fZsXOmaMLf
zVWvbozNFFKzgz1Z1+n39uTcQ9miPB9yuVd8h1qvW29//lkdKYrKL16Nfo7eZlMi
yUnM6cfVAqhxOmsgSpMd+Gp2EXQxSd8ubfT2NMjSq5lwcmsUAchFH+oCPcLKaICu
EfUquz7eNIFXDoYAIXwUYCiAP+ERrSy+8ayP1rJ/WKep+H1lSCAg6MpUr9Hy/hG0
7WM1yht3tcaMwIcH01ZFJZnkFyB8Qqkiw7C74aG3DolIN4wf2IVMUelE2IT8ZYHo
kTzCx7SGKkPjCeon2eTWreFwwvCdWO0GaoJnLL95fzmriIP9y7lJFN/Mv3L6rghc
W+l/0tu2I8bfJB6BwmRLzrW6K0vny8K4lajH1r5npZaVlgw/da5ZCVv2N4TmuhAy
2N6kWe6CQ33nZpgtJgGw9ZhYwcDfP4h0tavqBh6XCInh7qNfZk2CJC5b9KfAhpRw
rvT2KSM45GOz4bif6EaQd3dfOE8mXors7P6ZHAp6g9r8xTXuuOuUnPX9Q53ZffV4
Rp/liuPSUDmu0bZF1TzzLdEThKnptqmks6DiPtYfoJEHs+jTTM61ZDBB5rrQkIua
AFbuhmHIedjJ1J7sE/Xs2AWZ/7RdbqwmJE7M+b86FJKrblIvNWZGzXo2KRgXl5bI
sKNjza2IXy6tlNFDlcDic7+uLX58RsaAnKiDYO8K0wMRyD2N1h3Qbo88p5Tc9Ou9
8pzOhvTYtlK7DlQ64KZWdv9jl1+TsF+fnal+8xw8ZBWf+oFLWmC2nh1XNTxC5Mfb
IZafUVrgALx1hekYKxjEqgCf+p7qH/O1VD0axcy4sSAn88DXurnqRTXXuhNKXUc6
48n99FbfdyAAISdGx3Ll7I4hV00AUkabqEoC+c6BpvSBy9CvkLfZsDLRsEbmZjM9
pTiQtv3UdDq3sDHuPvQsV4cKJ9eT666Pr5JSj1a6eMzc8caRAqUas/HJys73avZC
ZqeTntC6Fr42SDPP+qWYrUhitcd9/6FuS8IUTGG58dntZHnnlpgtLb/Dm85Qtk/h
oXidxRTLyHTBsL0vgajNzTbNZTDFkNjtSNeQLA+nRwaKUnzs4Njfh7LT7kg8993h
4eIGjLyPZm3Yb6obpu2T2zaSG86dz8E9fkfnKlwyT9VjdiZ5IrKdlNHUOablOiNC
UuAdRZJN2GduuXqYkdZ5Yue8GffiBewGCKdlccDJdpb5aLqXGRB3VL1nNe7HZ3hV
4CtyBeqhXufAashuUkMNiEia82U15nQAOfQb/Ht+4n9seNKXFpJ+znXuXian7kpo
UosmA2Qyg+vPdl11aVtoLdJywu+sxwsTrMCdJA7TAyspDqShrnd2t4H4gDhiuuSa
A0lwurBFJjuEApVBOoQE9GmwbiTMQU9lVs2hpZSaYtXLZkTGtzbJWMUCEMVWtMT5
NG0232NBHYYvyNrHJDRXl0FcHQB+RzRIredvaO/8IZYCFKNRM7BCkvcmgjw495qg
YkGdeZeM2OTtNRvqUVEdZ2fdcwtqE8ul2jFDsvIQk86g96gC7WDoCHChmGO+FjYZ
hdt00e/3VAMa8jvVqfx9Y9nK/xTLbbQbDrNjJLWDpxOViG2S9/6+dzJV33+PXRrH
3fWsdmYIuxlu170c7o03uj3elDkzLd7ygLSmAq+3e4V9+4vqlwTGexbrIgOKH8jk
mODh9uPtoFzzxkBoJHSADdL7GdVptHos+CP9UlDV91n9jkWuMFc7qs6i+5AAopg+
6FW+rkA/epzFAhwlqxD9C8Ufud28IK/wQVgOrej9YZsNmkK59NhO51cOFQapVsMl
P1jbxUYyRsfPL/yROXumfKDbpG6tIOxgh8er10sVhhEfjhcBEjon6rPYB5A6Lg/5
3OOCaRTQs7CGxMZS8NAokM5yheF0smP4ZqzLDvW/8XyDrK0sgMV1nM4bDmKvafrx
iOYciXcAtvb/67sTswGWn3aKSX1kAhoAQxNJ8KgzZi7MUhNZVfyLjUrjptQNg0yv
3BTUmAveRdEvE7j2Gatwd76TxmzuGgaom0lHO+sKEhJ9U0CHnNPBa950b5ZGxWqX
Z8XxuW0vMsfJBpo5Kk1iTSEh7X60/kc87BNdJ5nBA0D0p/c/EpF5e+HPHMVMyrwJ
TSdUDTca/6ZsbrLb5+JPJ+FkS0uyVB9DoL554YXaYFVGBRypRzEeIP4YPAgBkFBw
b2rQwnMR09ftwMYKeiytslBOI1rP0i1wTFeU2Co0VfLiw98h8ti1Z6AOSGN5e7Td
gazhCkxtkG08srmwGtpmN53gc/SyCJLqXACyqT7DoJSRZXPWX2XQFaVDIjeob06y
1l4wE99tMkFeWqcyGEdnjPVN5svZuX3zmuJliB/N1tTicX3VspkBvUmBfBHU0OKb
eqg8uZB/lgWWOWPGUkdYSjyu3Typu9QEXKIfyGpW2EVoG2qbSHiSVYDqAHLikvWQ
vLMRef0X9t44qHVvIHJqsCfPqXyzNVhUuS5h6nzgQS4JJEiEc8tzTmruPmLzR3h7
6I9twC/j/IR0wC4RC67GzFnJIL8oJWBcLBpGAAlrULyw6iDhNwyGK/7RAo5LXBpE
YJULYUs5WyRRrGzuEQSBApmKcQj2CsqAUPgE+11VuAys+QPgcQ34mTz31xpYhmM/
exKPf2C5UrkbSK18Nl8w9XyhwaOu8yD7xGKOz2M2dMXVykkcWbFfmskRrAheMvSu
sizhpsqO0HOnNqj5UY5vgQeqeJn01o0pxBA0nyUVzRzOu/k2w8/J2LoLQRsASE0r
ufmTow2sOE4OrPuLFeo+x3zUwncSbcaX0QNObFRmvRjJD+6wc5dQQFImb+sgu6p4
1YyT1gF2vu7gUXuNgbby2yySQekjpzW4paGqAgHNCilT+Pg0BPv0TT+OZqqis2v0
M8XkfB+oJVQB8UCrfIJGVr3R+/7Hn7UR5NimiDV+YGhVC9aIKt6W+HQS2jymA9ed
6Ektny6D3mb7KqsgAOmsdoc3LaTNjJMhXTU6QmldH4VekrGGGSIxNucgrkPS10Hj
txFRS491gTRb+xMjELhCKqZGnPlzA7dxzUpCs0zGWRfKd3cPL1uK7WjA3COnr999
icDwUqT7Aezp5VxoUi5GQZWLziUBH+WG5yLaHM2jFOZ4fCTwT26yKIJ/HUNQsmGJ
mid4hoTbcOba3A6AD1crGNUVl6slJivjLLTVKp7ZurDmlizGMRYjIKGapCzifa4O
VBv3F6C1uMCtfZ56LrIwW7j9oOF5gG11jM1Q2e5Zj5x5aQveFnPq5qNiW1Khp89H
mBCz66NGu+UOYpw3U3ps0729d+yIkPjXI8qmZWMmGjyPm5dRlhzKbSH1UY/UYLw7
aHk6dLJL2ZzkfYPTuNKtFXhXn09rsq2pGm5OsPue++PfolZrMuxXQ4I/C2+B6ggr
agUhzRvjmG2BabdZz3yYauQMsGSKM3EuIZIdmdjTTSS48/X6oyuc+d5s4/HRD/kN
nYefTvoJ1Vo713sTKPWrOPGFPci+Wu4wKOgQL30hsYesmN3Et2JGW+xcC4mupRiE
cmo/36NdPGJUskF8KURz1FoUq1gARjN/q0QBoaC7o50dx4v++TPGYBBHBKNK8Xfr
2QayyE70Jf5+g24r2Jr2QhFZrzuNncidv3/PoSoryTNFANR98ZAPmsPbytUB9kCO
n1xFgDXfIm3N5WtoLoi+qefevYMeqeNXHivhR3XE8NL4O63/lGGkkzNw+nuhbSG8
p0aj3lk1TfodD+yGVAJqPG+iuWN7tdtlwUmZ+tHFwfyxo7uY6WTnulT7ObdOZwVI
GFEgljwvEns7ql3oNd2wFG6mU4ZhzxRc3pW5ZwNK7UThBMm7sYZZ/oanudBYKiEW
vuTfkX91nt1U3BewCskUSJakJLnof5FSEMns3Y3e//qQPdY+uvMUDgEZlR0mxggb
Sa5lYFc5MNjLNAusO4JAiitfYkJX4hnJEAujaYNDyvdFed7qQ464+lBs2Z8CLOt5
oS1YSWPR9bmwr77xd9wgy+svkjFS+a7kOk1oKqGffdxGXQwki4jONG4quuJK0LV6
TSi+jEkEh67UZn724A86ouJnyJR0wPy/YIrWaeqmFrfXLtCPv1LPHUW85WKBnaXz
JFI0VIcPO9j8z+6VSu788BbMYFYLWy/XQZ0I1YsmDKGYIsKwMhSw75w+NaCLlJWS
AOojxGGhTiOuQvfaWLaDm/JxW5aK21W6CvTSwDc1zUVO/KgFrR7B+1MTawZfTnti
iUl26gKc92VFgxFT6ryQfBhwcQ8o434LXt0Y6dnTsjcWy0IzLuFFQm4L6XsNvm+7
4bx0S+48j2SOHgMEuzBqnHrvSiuoj/RNZ9iCRmgWtno0UpD9ACOZ/87GaDo4i5AE
4ge0QnVtSr7zJRDidAAk2lgEfBa+UNNXfSRSTHkOU+19T7RAkMjb1tnzGWPrVqMO
wPhyZPAQBOFEkNbeY61Rn/izYMcrc9R3g34StM+E8jmWS8X2V/gTX7v+EYCyVUzR
sJ6g4YXHCXCLikzB7tPJ0f4eRVXMHAx6D/NrF5lP3bJOlJuxYX7ZzodYo6hK2/g4
kt/X4SsAPTnPfjh831FllDUDy6euB1Mhwn+PJVWYGghkqgBDuTVGV95TQBD2LvuB
jNCaQuJAEUYcTJljJP0AsYAnpybeo1ZftBQ7K3O6I2I5Bw0T9NTUF/T3cEc33YlA
sNmE4xVPt3+amcAtOfU2cP0tMySLopg86JBQSd45WKfgqTLRnQrllBOX9GviBcDz
qBw2MElK7jhPjxhG1Ijh/weIqjGKMlvqvPw0o1XQhQGEYmaVPqRabmLkQAJp6u26
c3Kul5iTlSVKFm3Hn37InL1MKlbv3ZIGQQco59ODDrARebeN9u309avSbmgH+0UV
ICyASCM+rTDJ1mc9JxWDcCwiTvZQTeNC3kb7efQNcynLrDM/pukFFY7Qa5yXDf4F
+knCNxQZFGoKwt10FPbtY4igOs2buQCyIztU4ldPHKPkXxTleI0a/lbE2kRgX+QC
XQmD0CpS4pvacILKOQ1pOYfCQm8CGbvwZP1Cer4K7d2+ta7ZPzWW+mIxjnDmfOEU
c3e4s2L84a+ruA5A3U9td42PHDF/B8HAPqJtieexCxM11nRIItdP8cD8QrjIFwd0
1xotAmr7RFQF4gTohLwGsYH4S060miYpUFE0ht8Ap3EEUrO4hcX+4npWjiXHfEWT
UHn+U2gmslYMJ2QgjRTYdGPk+67aYLNMY8DxH9iv/QI=
//pragma protect end_data_block
//pragma protect digest_block
8yOFcSKgilYfMlQb0xHjKNYEEIo=
//pragma protect end_digest_block
//pragma protect end_protected
