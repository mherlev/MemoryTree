// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:52 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
CaaQEZOidMbhH2hYa69GzP+bXqi8YOZ22AlTndyopvV13gn0EiMguBwudT5jB+Og
iKCKtVmUJm3C24QHAfi2XK0dSZWzI/YvYU49oaZDxqn98cq2QOijxwK6NfkuwouV
k3CvdYLgyhQDkxLGuua42SvmzEH+BvSgOISsmQOQZbc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9984)
dtikCcKk9k91xND/5t+HdJ2rSaAJC08O2HHmYmqQ1Yeib5AG1wW6UZQmai5PrEy7
xUIdJYM3xYuX2S1z/nSsLOEOEpiESj14yRCuaggWfrDBV+DrIGiHT2mEK1vG9h2O
S7wwFUL+pOxBOQPmXkvSMeH5k4+T6u0wnxxrK2EDhfnfTbDMOHpaylO0tGC9bj/A
TjPsYGUtQ5QrQaqHFHiiIYujIg0OTlTDRuTaJ14bTOeTQpfmm3Nz5ED+X3gDDwtv
RgzVTSJQGuiUwAlX3YR9LjJW5Cz/h9NfgNoE0oYkqalAp+FLAeetAYDHBXpXY0lb
sJuBFYQAXDIPVd0Lo3pgcCwnXefJtsJKLC1C2EpAf6xyI7cBJq3Qa8DtUCZBij5W
Td1+Hk4KfAunU7TRD3dS7LS1edIzxHboYS3+XSi9t3zKKjHh6hNkC22ZjFTtr4QQ
gLdq92QlWCedxanjjCGZwrvTd1GSRYl+SxX9FeocQQBhf3Baetm2l5llHz5E134W
svnmrlTasBc0uRm1ldaj+qULjGjqUK99YqPbcUUqt//BcHprZ758Kz+EvOa4lozc
/Pzio+aLnQ+eqexYfuW3t1Yo1CZNJ+goqkmctPImCLN9l7pP8efdWmBx5j/e3nmW
W8XagigGIQvDGeUm16DYhQhpAvl31uEDU57C/WTXhDAFjRJqWHIrGe2TrVSlFxpf
wy1MyxhTpPTPsFbR88Stc7N7cJafVaXb4bo7kuuE5RjwPGR9NTF38ulrUxm3lq/g
kuT6nHDhEloaalD7K5GJnQH+ola3lz6R3PZyll4HDRcEYc1MiSylF94asBw2llcH
S11RgbMOE8OXZvzSSPg4DVjStNGw3ysgBJ7HPTRzH9cY2kFDFkvS5kbKNKcz8uv/
BODKTSEn5tpvIvV+EFnC/+QS70mXdMhLhScr3VHDYke6opN8Tbwt95tUw+h2zV6m
+5OdafxaP8r+BhPT+rvvL+F8YFiaSDA7LRAPp+yMSRMiBE6rz02EkID6vajjHznv
eebOgyyp6TmF/21YE/iC2SVhVXwnZIsY/BJH8QrU7KhSNhT5C0+ElCLy8nO77C/0
L00lthGUeRe4e2z3nNGpEodwxeNnu/EjLpG0HU0PxXlcvEh63XurNQxyrrXWTV7y
h4aHqRjObLpGlkuUeC0ifHWDwdCpP8r3hubDU311O5TZ4yKjoMiu9rdLkaccMydh
Vk+l/LeRPcZYX7Bwqu51GyjcKlYQRzDCFVjUOifyFt09dE33xnc+sPidPV2DJnqz
NNb96xJOK0Se2n/fOtDyOWoF54+2qLOmLgc8uJxMMsJj9F3gRYidWipih2qta39o
I0TsztnlGhXCIrr2NrB+nZ6cIoeSOo0teFNeyjDdtFwGcRm8w4tutcG4iejILA+M
iMsN7uWKmD5kEat8wVIlJM5j2qyjQvnlQxoUZ7gz3OMkKJDP6i7ZDL4Ugoz5tmoW
a0+cu42Q1soI+zC3byKk2GnHat/2Y4cAXuUgWdjBBwgS095ZgLXbJiUBUKAmFoTI
JRARd1Kf3uZ/SOkXKQQRlNt031zDhBN66Jyjw5KI7J+l07VkTRnySkt2LgeX/OoP
nZ7pXTJxxEWkLX6vKfXRdj/fwITMJ58odCBnV7U+vgn0nMqOX8KptfCYSOFWytDN
PGGSySeLNz/ltBxpRsHtMypUGbgDsRV7RmMjZTDzNPfesXOJwyIkQfHNQEDmL7Ly
KYDKTAl4u9DlBbxEBEDmZVgdV0agJAxXlFbSA3ahhZ/sqDb4ivOWeF9K8M/P/aPK
vP9YWnuoDmIhnXTzl1yLwmvFGFzrIc4RULsX2ed/NYfSm6ub+xlXdMovSZnUh2S5
WWAlgp8v2nJWvunYLs39wY34xO+soFrPucRw3JBzR81GAnTJhIzfCGLdMgk3q2Yr
RZijCp9TRd+jSDVIb1YXiFygMQIPic99IYungNkXL2RbEfRL1JW72jGrWSbXk//O
KazJKqKmvcmir2CW2qc4UwdbNmhGnda3BwsDBbtynTv0Nia0HtcyMOMwyt6pBIcT
CLbhxx44z8+Rxe+GnkwE5tn6sdHLtOmao7RIQywnhmLDE2BPZN7zeHTYr8fzIzOL
s2ThDMz3qI3BiktCuiVqvC5VrRJobgLsoawmxyBJBEewZQK8O+y2oIwallbc9jw+
2JPsJcxssGZYpUr/Livk0zJ/+3ixqb4HPoFQg0C8ql/PWKIcyzoMnYDBP4xUiMGg
GGKoPtk/69OTilS+MNN89LmBpH/jf46tmZHhc+8zEUzDdKvRSz2ij8fGicoXw1px
jm4TijYORimNdtBwTJ8nfO8gwDHqHrNbwiQ+E1haJBcKHK6uhjdKaWRJkklZhxc3
VZw6A40BxHcVgbalDj4kGPBr7pt848cesWhHJHXnEjs/qnROqD4mWQ8w84THfl82
lauWv2VgZr1tD0sjMkq2OgC5XTRiVYZWGmHRdX+YktfNUoc7RttH80nMd74qBxoP
7inPl7/0mO0oIl0vydX7YlS8nZG1YMGs7puQkD+XEk+M+8wABZKWOFvukENGhZcW
G/AZKKEKTW+yFqzZcEol+NiaUPQNzcyr5jq8cN95ItrhJkOQ7HYnTBD+uWBRJzfC
kRBGP/a6Rxq4kPdC2SIUutIrayuekeftIDr1InRIOpB7klXTuw9nmBYcugkqKwA2
Z7fKAtnNxqXQv7vDdwxt83L5WAOXYA/Lcyuk6yOnZ/dU8sPdm3DuWIRxxFXDJHrR
eHNfJnXpNGZxwLAaOcpawc1Nf/e19YTAzDi5ujIV9J6BV/JyTRqhJHR3xN+DX1ro
7igFPvbO/Ab+1okvDX6ua0jZf76VWe/2eUZfZHm8NIOMaZUJUjXHEQe+OHfg/ynl
m86b4NRQO1EnxDL/kxsi3xBaMzv8Mc8xoprBiJ1M1YWgbBDvIsYL/lfSJ0tUmblc
fQYQbJCfmL2ztJbEO02Mm7+aFFuOHpUdXPx1owl61FZ6e7mGkt7W020g4T3VpsWX
kCH+xbr9r78blwEumYCnVk7AUysuAAFJmrrhLXbIAnvQ2ibqSQsGkx7mxpTJJrHX
a8uZzcvkY78uu4OuszRFRfhMIHX1HZMxvOCgkwy/2U5kAEFZcbTETCe4+kWy5m3J
TTjZgL+jq/ce/ep3YnD+utTs6+xgGCmYOEUBXyvFwRYT4Ng0VdxEjmPcrSYTX341
FKICexo92EN1fUPernyq6VNXq4sF/M0pJg0uQbObGXQ+DSr4YCrgufNnSQssym4+
exWWDpYOzwqrNPCy5lr9aPEYSY6ROZeNMUu06IpUIFGgxnKE49duzvaR+eb9+4V9
6Nf+QVaYKhsPpry3SRvV+cC7K4eI+M2SRJhYQgTQcZ0+qwtwrHJMXJYenYu07v4u
O77C9pNphDNzb/p6pR2VlD/4n7kXxE1PDG0VglXzN3s0AeulANnTgwreD8g7IIEA
0HNM8K8nps0rqgo1BPnZuNGDN8jHtA1btDJMqG3nAjs9V9y4/03rZXDjKnoDomEq
hv3F9wHtaG5FRZoh9xxTL920NUvHaTHGKuixrt10Yms/PrBdOINCUl7eVlxVtQ40
CKLI29wsLOSzO2vPhFNYcgCqfZa1y8VVVNmgZjNgqNlJaOiOQfHaAI2Re7SbOC67
LrnbeRuoxmHidcjOJbHVGYPCtqYb5CNd23/7h+mEDU0Y2LsjoMortaCZwR1/8ZDL
hemFoCfcKkQRbIdlmGJdrFJ8pseBE5YKy65R+nkPfeaDPDdmVZH3D8LfsUAhvdYS
qqDctEDx/KAcffxHrc+odIeTBrl0+wKZxBxcZTzLnyMQdHTdbVrn6LlSjaMsLM8x
CnJmfPKjJG0I8U2QISjslGvbJwwzAlG47EFq1WAPj3DGEcXmRP4BQBq5UVCIU1In
nsc31qxkN3leCpzyXPf8+5V87KtrAhB3cLkoYMKBV5QZ7ulF4NoE1+4TsTNnoH61
njxtBEP5h+ifbpqds9X9QyhsNpcVcdMkPLHjlNmdQlNm6+01qJRqTJuQM3vEACKh
/aRfjhBstTtC03b5I2LmtAkK+JeP20SbR2cfHQQnAU8brSPvE+c1ec0Gh5cEC/Cn
zp9piqwJGrc5JUXOKfKeoLXPus0jLt2xFQU4wTs4IgOBq+10KDVHim2/ribMYy1E
JiVtwggsjuEboZOrboTdM8/Jw4SIZsFhBesGnwDeM7FTNnw2J9v61IhY+o2e7QNW
03LJYayydUalxh5VND83DYKC4ng2VAzsdemBAJnjuDnipeMOoDTvuHYblo+jQyhH
VqH6ibh1jPnUsJekTe5Oxha84yTTjAHVzt6FN6LWN7/T9YHrUakjn8sxfCkAI3ZM
iXBRuRDpkK2Ig8z5/LwQHR8d9InpahahlrmR9HcoTeFz3EJGMbNTz6Gq2xAmIt7D
o03iJyVfCROIEdFLBm35g2LV5rpXniH4IZ+L/hfX986NZLGqNza92NBP9k9CC4LO
iG3jMFsJ7I3Wfi4vsFZKPHbPVBnQeHVgyFqz+D/UMP2ahIFnYIj+yg197VcR5dbS
CrDUL2B3pt6leTeHAQFSTjuLG94lVGfuLwYBeXs2jjYowyE6MHpUpiIdMAaKwceB
BgJiajxYJQ00hiyAfOZxprhorRi8pTPhtayJo4u2qIfAjYUCpNj9khc5IcYAEErw
ciYfuME+DZiRzRBML/v9F+/e86RUQi92LKojiQRh17DtEG/EG5D+3mZMYQX268uQ
PYZ5mRnl9gSJS7jl6KsUX6Ly3UqThKoBBUaA5L/a1xKNuRKGnooFGlhOLEBV+ndY
0YM1WCJNj1NhszB7pWDkE/7ROkQicVoxWVA56/4AsjfQPY8DMhthiWCilsF3sYkl
ax2GqJTVKYfsbmKQ+CR3uH45E/mCvKhfDkSOoLEiGeZOz0u2Cn7sGapqUgGw2HzV
FkhGJXkP+ogEBJeqa6/IM9KET03SvHmEooMWTE9fXp6wy+E8czTmWqxd71/UAEyn
yG6SJCY9EQNwc45rD8mHEDGV5rkpD83W5HDRm2OvzLEZH3LTjMnusknUujGwUjMK
0rku21uEHE5Ij8mTSiWNh3t+bvcoCZOkAPORvmYtfAcULgbUtNDqmWz5vtqByZuR
AD6N6vKPciL2/HXR7AwcNSww8s9zNKMT9N0iUo+Ix4TEFv/Oabd1nMJ/Z9B8tx2N
yAWnMIsGJGi3CPPOd+fEkVENcWYbnv3fL/WmI8TN3OVKLNrYgb1ghv8oTaGOGFYy
Fl47WwkMcs7Ha0DaJte+9Q+t+Q3zGJEOn7lkxp0w85btGb3kG7ikPU/SW4omXOAV
lNKsI3sUiybDAJdgWvyMnidbF427WY+0BkUo4U9UPrazWyNV2tke/JbwwZZcFDGl
6fIyw6n4zt+MyP939Nt2LvD6rgpJuUJvVPXDhDGXIa8XFp6rVBCpdHtvD4iAciZ/
63fSy54hp0eJdzQfQkCQT8l+J6o5JqQC6IMwJC1lPP+tgvUsXXGleyHpiA/g40wX
TMAIGUDoT8EDctIfadMcEr1iE/oXyiojfoj24+pVWwpk8OvsMFs+SX56D/zSPCFu
ThkpjIQuL4NZvZBn0I5f2reyvt2vHppAKAFvy0lAtQw0BXMdasiumemouV+1LLh0
x6k1SAaThpH3aCAK1NJBZ5Xo6VVHHX/6xD7d86o17OTWkW+X/DBK+2HNhpvVIFLg
7juh5FBoGUM4Xsk3kmNIuBdi12F2z4p1kktq1dYxULD3ow4BH5KUZFkqf9ptTB+N
gFAIhkC3HW4ia/t7oDmHN9CxdmX8NE26b1NyWOEEsrOOzY10hwQ0+tfaC4ay022C
OXtTj5q9nVcpeSibUUjbtWcU3/ey/w5gILZuK7qBQxKjYDHilU9tfpJqJ5Xd6VWw
bVa3mXwiU0BHUcdZMO/d0loa0Dah/JR87ZUxBtootgQPZbWtm/OhS8ZILvRtnIhJ
GcxLYhWc99oEagSc6gpenQEIkDUkurww6ULW+QYdSN8CHKM3kBk1MlmiqMriz4sA
0ddYF9HvzLT0NGJ01K1rxsCQf7w27XjsJjVQ+s3Mwm2Fa8Wumn2XuO6fs/kXrPn1
6gyFPe5ObJalkgUbCOPKmS1puCVcG1u6Urplk/vhHoBBxNmHniL2gjGgqCerkmSE
Xv+zg/dg2M/wfSEq3DrTYAMBaApPJ/4hy6hbLU2QL0r2fCu/h2fAoAD9+F/hQzbu
5HbrGLFSfvUAq3FcGe4AcyYdFUhj2PA1xc1q7Bt7krJm/dTcfLflL9AT00ynJLEX
d/MoG0IAj+m5XjF/1L441bVfoWNoyMAQh+L6FqDgUeAGefd+oILtft96mmdYEPRB
v0E0GTRzJBNtmFWTytseM3lS7Yqq05IMrSN6dH8T59iQsanW1b8nrdmGghAXiJPV
H6n14AW9ffDrgO7mlja2PToTn7b8olg9livQGna3Rg/T+pbf+YJBRLDtzb+nMfwl
GxsJVSSpgnGJWa0Lrr8JwkrVOblOwj2hzdvmmKft2+c6QJV/56gEj355FAucajcT
d/EetAUJ54C2EBjV438o24tSzXdNNp1sAhccb7sYK34E2aT45ayCXwVcsL7Ijzs3
pQ1Yhh+kPUOyw+6JHV1hbr8k42JPmohWdUhMpRt5C+7/WGvDasHuHiQMk5r3/WNH
Bk8FcRYGZ7Mhvi9ap6hw+AFIzQb5kYw+NFumfuLqhWRoLx50llu0Zl26TSon5Cyz
BfSJv7wWRDVhxw/t/WIN666Kx7szdt9xgpyahmx/xzQJsHWVxssp9GMOmlikSiG4
CBLLJgqAWbGq7DeP7Pf0VjNaUalafbXO1q9u1r9beedxL1ZCsjpJVoYD473ZSSDA
1h9sRORVNNt7WOTRF9SJrxUDoGChdriJKy3SyuEAVbIIzo22HRajsXH8SyoIYwAd
JF7h+cvWitFJYiAoUyIZz4eiSQk80vGV72pZjLfYrYkIZADVr1KtYk+u6c/KZhfA
p+MAvGpOnpLu4GeRR5SkOGe2y6g6hXlE8f0b0lwfeHKg/+84b03WhI8auTnAK2ZR
f/r9n4w7ugAFBgMdPVGkCSpFHFABuS0ztLdJCH0qTPqAELcMe8Kpj7tITIKSdnKB
/bN+vVLDSyA8kTRzDJadGSLRvcUaA6azvQ0O6ujeyUMEe/JnZbBZbtjOJiaumZC5
v1v3n6Qk8jJW3wuxKt2lakEF0BKV3neos/y1l0g7AgN7iP/z7R500pWVjxC86SRu
S+aDNeRXwUIHdfl1X4oR16HG5EtpdYFz6s5jyHLSsT9b2xsoilK8XnuHx+fl6c9j
zEDRIg+aLgLaLwrn4ekemORrW/24WXwXjM13QdWhqvNz+p7N87pmNBsUPBFLVN87
2iJZdrXTndBuG5dGzugUr312bD/SL7ckZ5DrdOg9KJwOz+90P9mPQwUy2yiGQMIG
rOAxOdnx1aymjBf7rBGDt0hTQFanElmwS67wOyJs2WZaY1r04Pe4zwqoP89wQw6u
ePCq6X+NVCSouA/FkDq9En3Sdc85k8pE2yodEx1F/CyWY9CSmQMcHUIH4saSMbVo
69FJKFsZJa9Wfi4xsGnrJyUl8HDnZ50HdALr5EsK6nenFIWIlQDObsktGBZVKQRx
d5PvJIrDpzUbIyw5pGjnjlYEoVUZYZAQEAI0YnnhuXX4dp5Ad6nYOM00xpamkiMk
XoQ1cMzUnG2N5jANHjd9JKW5xM/kdw25WsmgaCrRWJidq7IwsHwij8ZP0b0zudgY
/hLWfmF+vBpH7v1OaI2Na/XQluaVUe7jH9i8pMM1eL3OOP7UrvPxPjQMkguqGBrI
vq4U8TnOzssZBINfJArOsCQAs6VkNnj7tm06RjfVBg9UhYdT30bS0kBWQP/gdJ2h
qD7/D1u6aYKSW6o9TLH2WbW2u+p9+zgq/V9AlvqY/zIqlxmLZNnYvYTvXOZH7qbB
SyzUonZeiRMIEKjb5VBFTRzOHwLlr5uYa37LXlCHytNTFRAbpvMiSrEz0jXok/l5
7BbgxN1ZdY8oHq4PBuybSjKL1RpZPO7R8xypOUhNStS9J/QjCjdBb6ahb6fLWJoW
SgGeq6axlBI1WukMlwN03A+I4EjJsEWBNwfeEmUPp4+eZV3YRZ/2Lu9HHpIevR4/
mrklyOYtmQVvRuWxflzDm+z4zJvdEo1oEkvjCp6J++tcKM7qPMnoGPGhNgazeVbP
TP8vM9otB9Nu0ZfGvBC74NAS7vjB3mBeLQWNlJkefS8Sc9TK5vuSM32m8oHR1Ayg
6bpQSmmrPOTsPknaMvSRuR5kdrDQfPfUQYmzN+QWuvjxWQGIXEQ8pqca6EYHVkEM
PSZOGoM4eR9BPbtUL/vEBckjLTP5n6N8MKXK2qK/aCuTeUPL1BExzM3DjFkpcyhH
i9S9LuD8KpZoz6XXHBvSwKVJxAR/R4oW0VmDb0svEiF6VgA2mtQ9lgqkJ+y9Newc
CvBb9RIhn1Sp87Oana/mW+Vr7uLioxkGWH4XN4c+WYx/Ub0nr0RXb8KVPghUiMnG
6hqEOefZBZc6uBVopzXatbf1RHnSpbaL8wyto3Owwi2sjfCTAuG+ezJnXVeXxyYW
l3YJiwEdcE4thr5WclZ5mWtDcykHycpneXdRwnkDqUqd0FMO0mkhMOqqjXKFsxv/
nd5qNdrnmJQZzzDKuRXGONTg6lWmIS5+6aHp6HuHEtf2MYSpXi0zM8KfRnv1wDvI
AfDNqEFzBGgEwVdsEKHqbjiOyNLOBgjCEFCSC3Kk9FUe9BfcRq+UNK+eLRLhU0i1
BgEplW9LBinv3sUIsBJsgfJN8vn+kKiQpx9bU8bChcUYvCQGzA7nsaLFTid0WLIq
yvl4DVpOhoSYN6QnbFusZGAYlYrTJ9Przr0UPbzEhck1aS2t/Pv3AeeMdSsNYXyz
yOqM7yjXwq7mn1vxd/fVdyjfgruABs3IX0LfxNJTJaXy5zxf4/nWw6txc5jmiP7C
9nGoeKjE42wcVUup0qlFcqlo5HYrZA07HexKtl9xYQ5y+7pScKkXePYR8m+r3wtZ
YcGc6ZirQesQ4LZsA8keAQMs/Lzt2AGrIK5viPvOFXkMyS/fdi2uhF2A3y46Fiaq
f1CAuTjjG1EtyXf6EQJjToSDdxgqctfdCRwI8qlCz+wj80xATLfwMdPDl2AT2tpP
ILmu9SP7/GLfJdqS4ZNWRhyTFDx9iLkA6o5nsBmRVMbNyPMqUTK9MF0XQngez9a4
o22Gvo75yFmyFNLIvzGOfhBg8d3ukikHHIfQ8RYR8tYwDRTea/nBsW1zlZ2cHRFQ
X/Rif6225BErFW1CDklKgBbrsXqiLho8clF3Q+JsrhksyXuVJkIiwYFwSGBJ7rkG
N/3+dacnjawNqYqSFgp/dT48PG3gg/i0WmqEsm/3YVXjdPkrSUwxKdcZhc66mzMe
NjO/ef5t4mBIVn2Ny6cJ1yAK3qkoPiHbOHGMeU9M0E7cozBwKEkDdgjI4OyacAGo
tbkrOn+SF288X3a+SwXJFxv06i/i+CKQTFUnamZ2YsGQT+LCtXiKky7uv5XOgwxc
fn4mIh/Xq3CDGFl4bzGbJY3P1hMlyucG70eWzBtO+3B3K3jFiz7q83g/OkNQ5VVK
LRkwnKI5pNf2Lj8XxoZ6m6f2/AbfmR68H/kSz0GMlGM0lFc9j7/j0hFGEGlysEag
v+UdJNDg+YvXKZxCrJFUbgbgo2SgQ7x8Ahvk6GxijvpOgwB5oOy124qnl2uAwvDE
IvIq0yIuTG5Zy5ylbaozfHtuus2vyEGESFIHNXXxkhF0NbTFyGrm7mosmm4dNBm0
q6wr1GO4ahbs6/564/PVuD93F3iGE9WmVe+fIZ+B5Ff0/TjPttY15OJKeEW/8X5Z
c+569yNxR20RpvG3iL+ayXv7+eC5DAWRbLrgj75vd0G4t03wwD6ZwMX5baFge75O
LzEGVvY2y0fksn8BSUK8VjypTm+kUPt9pklRprXVfQNoa/rIZbh32njw0eETEO+x
ckzCrGlchMb6DFrPDyfd69bCDVxkWGDqgf4g2lTKO76UKTIUhvc7I5UA7gv/uYry
BVNaE8ZteekVLBzxMk9jauPSH5hGitBGMrQxMrV5quHC+/j3qF8/fpt8g6bpmnFQ
pVBJOoaqDOfkuBrJMQMiC4Bd/UhO9Y1aHADjM7WsV5mrMoAK1r16J3Vyg1vk14Re
+I5wnDHBMvp24s+aZ+aeFqG/owsoBzrCzxJiEzJvAXGjQd6JZFO2ZRX8G0zGPcA0
gyd+uD4HUd60c8yie6LfxtMapUwXnwnNMCcnPNVEWAmr8ZaV0amRAhxHs7LHTvrx
UAziiVios06IeNRv1GN7tm5S9IYA+j8QeGMzuCTHkiibszp+jeEToSUxU4R0E6Hk
ER35AxxWqaLeL1swCSvo8f2D7Y1RWQP8oanx+lsA0U+ukRZMCBHMvwLuwJg/BwLQ
8zF8NSM+Di3LsNwMM59q6It4+uOWClnL0HB0gs9cyXHG5Gw94hRn3ejrx2ioIFNc
FYqp+8kekhjFtW6N14gBgnoaCIn0VntYu/5Mq31InNszQ4Z2a8XAQ/cB0wRTd0Y6
ldfpb5mdJEgOoaNxtm/EMqRjCdQs52tHihxSoB4Hsj9M1lMKAnHfOeaBEIhRO41R
9ZJwXF469KDOuOZJE6+3mkV3pLePtU3pGgTTnlKwTmfi+/xIgAUm7xztYPclZwtZ
13QZT55vTidU9+KPI/QR+PMeGNyyc5bnwPYsrxZZvwntogiQnRyMU+QnFvR7/aT0
GvCuY7goM3chM0RZpK0/VQ5dMaBXS+7UbWLzp2kkYqIM2PhBHoRJzUHbMFSeiIfg
rdSdLaNfTYXv4Z8f4dhX7HVaW35MadFnQtb0nFJ2+WUvysS5mrh/en/GYLjc/aD5
sXzVOtZDrdT5dv1vmnMWJrgtYuxlsa5AMvKEEIlZtx56tVsksFQGSXxVh1U0ehvz
yv2CM/zBI0i5wjz9Usd6P3Hd9lGaQ/rrIc7mhRc8aU/sDHVJftiTuQJZx/2sMYNV
Ch5XftWmJ9KRK1MwI5+KeJPnhvxTq2Da6RzAD7nMCWRXauqb2i9aJK9esR9o36ou
JK0lU4OaRS6tWzlGrPqD+w4rQQW4wjmXCdRF55kfHl9SdANbUlolyRE12BrqpRar
2CPElItDOk9xzYyKXefmokNj61PGMZT/sdKWg+sALJE9CnG2m1RD3k0LPQFY09MV
I87H7478QwtwFdPLBU6UE5BTyJ7YiTxRinO48EOXVx4ZPJLvHKkR3H7KfaUHD1+P
Ku1KG3wiXh/86YVrCcpYb3XbKH+DisA1/OoCXm6/fxdTEnSPQ0yrfQPYGJB+2ah6
Mz5zMxxuB04tXwMxdRR6qhpJreI4yeBG0hN9w7/KVmCytUUsCTYLFKc0R0e8Qo+b
MQ31a25BN9V1IqFkY07lBCaaFaG8gAmmU9htaIhyt5xnMBV5nBSG56HqewW/i1ZH
hbCUD6xq5eprZB/g67vL51D/CiGWCfJCjm85GrpPYvNXmuWQnKoMmOh63CHrdfNt
8vUdznZdLxl3nsM3PcuThcqtLi8VzsHFtzBTZF80a0724H5c4j76Q1RgEg6gIiTJ
IERTbwl7aAPD8oPc24q4VahQIOmccXT+r/0ZQXCQjn6v/pi5by/laowGh248tl3E
x47ORbnPJq7/GnRzIszhBuWF7Pqb+bqfi8z8E/DwInQmCb05XU0BuKobi7ViGhkJ
hFVLj6g2gSKZJ+zo/MlbCuI6lIMal2GAVMarb66K1rbRyJPb7ZZAiVS+LIrUUKTR
qBz7lhURmGEcgW5I9G8rRK+Nh1SIOquLFvk9Cvxj5RzQz3IyNLsxmXJyUmGfTpXl
/kqbp4kS5XlWyCRi4aPL2BqNEvIYm19iHHp1rFjXh02n+iAeifgpisGvio4yBVq6
BZd6ckXKBFp3pErMTDW9V2LYihb2yduzwMCjlY/nnNhPwZgyTP1agceLkfanGezr
KU1TkgdJYEchqm7SxWLcrjmviMx2dBSa+sTlww0Ott0DRkOzzGttUeDBYN21ngKQ
WqpB+jWieUauL5lTqNpe2b5xfC+U8dDbVFwcXwk1YFm32uA7tOFRNdhke51YgLC3
9BU3s15pnkRXxg+zZH6mXWsWpCnV4tg5MEsiaXDxrS12BqD/2JLq+C0Ie1KVtkmi
5EptEabGTH7It8gvGafhHKZlLcAxsNfRqmXiEPTjylMBivpqKJfc/Cd9kOkj6Zn+
PyTy7Lm9kqymOTPp6mMS7Tso+wC/nw35hgwyPVBe0Wo0Btfnr7dQgCMqpwVpjzgP
bUqfgSw0KNCnRk8tZgrK5klgvgGGPODZfgYp9Fiw9mGNCZarGsb91K3ZEvZNieb4
hHH8O5RuTSXoKIbhe0LdWze712PXHNcwBcPkdkQmBBhOIFz/D/tnZtxsidf+bH8E
kSoAjr64gWRqirRxAK4WPQCUnXHs40boGQtGmcdEYfohrm8QjNkQ2QghpE651RgT
l31lAhWlD03/gvK6wRy0KUL0RwMrYMYKQq3mA68cJlWmeIiTqMhMQ+++pKP7mmgE
mvIOcrYboLvLThhU0J4c/LxXDDUksurUiAszpwpxC94s1AzD7HKew2m2+IKduoOs
aMwym6qSJ7G0ywosRr7lkyjjDvoUY14kAINIpQVSRoQWm3SKRXaLIGSoLruLkxOC
kpB8mQQRltGiD297fmoZ/G2c6VPxAnmwFvsBAqFKy1RkTCQm2L6mz+Rsmwn3LALF
/s63FwToRzwyF42RN05HejMvJtYvDLCTrS85GsM48k7Zd6OsmdVS7mWepXt0ntK6
gpeyAKMzLXXN1iS/QnhJ0efnNBTmuXowzRcOhcnHqEetuT5VDqoD07cM5FTXBKrV
4IRnooV5Sd6tNq2faHFa835LVrBnw4YaX5JbjUHrMu4vov1WvL01KWy0IeYlmbP3
aF2CnJbIZqOwqjF8eEuxLESsam2uzbSotkV52o8lF83DcJwrGb2pL3gIWmEZIxVc
s4rnhGTmnXKF+4bK1TngjWYrTOc1/gTpCHpQPNHN6xqexSUqJScLtUp0CwBjCj4A
MOoiua+jtWd8sKTm8ZMt09KNygmR61GRMJshgIlZZV34ZF5Ia6IiytYqwt7yi0XV
7lLkmPAjHU+FqTLf2vCvcGuYCLdqm3roNo1Nnty2ovtYcAXwReUqB9wFeVY7+szW
BXpBycsry0I7sJTwKhwZNRYiS3G24tW3+PYgmIOH4xWRSRpF8rQjFPvXOLTU/bxB
C0iXsQty8c3CONhrU5djJaPUwW294IG5i9h+kOz5S1SN10ZHJuZCZK7RKcAU1Nmt
`pragma protect end_protected
