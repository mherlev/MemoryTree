// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:52 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
tSRemlwEpBmkYRbKKaEeHVHka33e5ot6IKX4IrprlBDZK/5G7MYXe2xqV5p0wYnI
EIZaDDkHE28dBohZuUMqgbAKs7V9f8qL8KhoxumN28n3WOvSJxO60wuTBVo/pSir
LT59GF6b3id7ft093z+OffelIxAfD5oWYUXOpD8nKvc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6976)
EiAiEPXUkVmKOlQMMscxtapUkGlSmmZs1dYDY8XuuoDKcMVuYqNmDIk6WDe4DTF3
/52EEv21a7+8eInwxofQPAS8Gw99hTnC38jH5ui8H92/osC+kE1cHsdIn/o3mF+A
mb57XB1oXevfx3itGTKVN5SgS60NMO+La2kIKuHb6wplLqe22+aJcVmxcWpw5Lv8
+eJcStkGyk4gKFfqwpSmA5+Fmji5OvoHm1T55p2WfrG6TFX5cor/EETLHyPOum55
d+Vk4sQ0fs/5PY0ebc6Wxf4Tf7jv0PPy6x3aG60RR5qo/k8itGtyE7B6rM+qELjO
EGLd2WMc4fJIsKiu7xiAvOEuu/Ku3oxw/x4deDt1h8VV5QHaMO0yB1xjzO3FWKBf
Jyx2r+uaPhyeNyTVJ1AD7LEmXGKvW0U9ON84ZGOhkXFXcLbLd6z5aLwlr5qLPojo
gUHEiocsRa3DMh6mMB3O1huk11zcBZhx6j6aA8841bxh9UE51K7Q8zS1cZS9LH+K
99zGrgDnGU8egbELCCzNngGn0LdNOnrEPEzefUdw1ZEr83RHk9exyIFFEJ5BQn2T
KLV2Rrs7Hljc64t0GnI5KXoc/87ToqUHTxLWZza7lUHNqMgvpW7E26CQNGH8ccMw
cm670RlLtKOtRK9YE+elnkxeGDRX3gRyTsPMrhR0RbIy1qQkx9sbsEBdKS6vO2Bd
YpFzJr8kuRkpfOhDOP0JsH073nRE6rZgOKoxRU8ZHSAkVez37igkr+3dlPmvkz/p
N2qPSV2yRXFy4gsOoQHRahiGQkKY47E06gx6FidiIYqdtBme6q61s1I/Fniqudoe
QXSgN0Nzk10cCjG65GH53OI/eU4MDWDDR0rq1k/QOdMxfIlvcMkXsfKY4UX7rhME
mKG268QdcshOv5IjPBMPHxdRWybTp196aK/6/e8FjiA4aZ/5Sw+ld8lOGCg7A64I
PRlQlA1485aACDjUieVY2FaZ29iixpRruqCg+Y6ggfxC3tdJPWsoetSve48yx3H+
QsgSN0RFZv7LtskkF0ExGr5JzUR05AAwgknfGKomO/sMLFAkxvSUvd/mQNl5vt2y
ILC9Py4/IVozsDnbSrYiV38xe8Mrp91Xah/txWxzWYOJe6GVb8CWwPirqGWXcrlm
34sLkGJYki3tmnCYuGYl1iRu1oVTH3o2pniOAxpqxLJnXoFPBVxFiE/7fXY38XaE
lvLB3mNz+rAXCe5viDOJs7n0+LH3ytK62Nd8ZyAY/suZFfnUXpzOIg2fi9v30z93
IRcyZiJIyS0dU/DD0bZmUnIjjNt56h1xTojoNsrGuRkbTNPvpkuvbyfBONqTMr3p
Hkuhl+L5eTn5exoCLjKmz+SgpQxO0nY5A7AQ/027SkuU7TaLxFbt6oEadjae56RA
FFI9jhylPBkDiiytmmvFjJopwxBqroW97wbcysuUV/XI3rqpWQNCfIGyM26/QtMn
JCFCmlS0qHbtgBbOXLZwy4B4AfMSmj8YN52mKEXlfnkpAKj7z3QC+/ivWrY29SMH
0AU1B47GBapMVAEEFoQ2HnpmJoWTEZIRX4qMcVy2xRJ2pks0CPH6TVaUBLHTByUy
DX+wv9GiLugDSB74W9WKuWdV4N6zZvKKJqsH/KcasCG8eZE1e7nNHvUEA8XPDEJQ
7kBWOwiUJoACWY8bdy480vOD3nxpUgWUwVN2tb/K4ZI40FZf1icxYg/iL8uPjidl
0X90A+nXFSurefPSTyKU64EmY5u4LO77n/WhRgrNE+lbaPHsA/2AnLYlQaifE59z
PK2Hn1A9mLWe4Z0yry1vpricWjuVopFk/JH602T5k1nOZ2GuC8HPzzf8rkRM+5JB
7rRmSQAgbBx0nsdN8TnqnNVmvME2aPX9bdlepCyvEaV4kPQvZah4ewIztIvBZuLC
xR5AS5XbtoXb7CMXDBkgMZn8QVzgniAwrIYqqELWYlAVfp9mJ6zdYzHShhsrHQ8Z
I5YxvXOn0ufKJfK278J0GZ1KjEXaJXX/hEPneqSpXW4jZPgwohptn5BKf7JsIWch
DlwQW1d3zt3VZMUaALoTxlTR9xocC8IchM9AmxoRbrRWCubPQM5ZkKaqPFAekvPX
eLBqVYPGBdhBfq/hn5bvLjfzubOPJE2pPjRIGHKHnq+3At/R316/ngHQAUwMXZDn
OGQYxPlweG2IfOt6pZmGEUbHRXF2E37KEYztQE9R3E7pkAdl9y6kd4Xx7U12zwTY
jvIbQDfFnLK5Tm2Xxjs50PofWtgnRoU7Et2tVjw+XhuSkZa7FzubO0CRzawA6Ct3
b3Jth/DYQJjM2qO2n8RC7MO9TVl2WMaJycIRun260UqtxQbckr5f3Y5dEpxAq5RX
hDKza0X4WDjVWkgar+XuNTKRy99KAuu/DheU52MLfCfwGlu/lQBndbn48712ZjLz
ayvhcw3DfXfNZCH82oKmMQfNFuI2C4nHsqV4hZuPqZXxJXKKHVjGeiuoQ+pfx9LC
tB7eAeh+lDOG+a+Mb8WEl7UkPXVsLbqQ3VYXhVJEJudvFjt5jB6hT63UnCng03G4
z5KEOM/jHw4wTcHXLFYW8ERmiRelG6BQqf+290Ad1NUo4B/yGqnyWIM1E9BLSEqk
/Bvg4OvT6KKf29gYUT02l47X2Wyo8yFJicpZZj+2JKrGhpKLZ/pgTj5OJqpP9L+x
kILOu7xCvtOCbdRUbgISeKHKCxoHc1cOJDQd2ue2vo1MXVRk1rTjSU4IaSTTdp1A
rWbMQyMV6ugGkO6M3DUsXPJeWUGGiQdalKoucVjFnqQ0z0yaZmBCpQr9hbzPAf0Z
Yh266z4UotdASszAK5dOik6rfl/RWo9bT4F2S3Df18CeK8JsPJefZjtI0aU9SOLo
5Jvs4QXn3ufkgqjpcketFe/WJdsGOp531vifH2UH5xXuzyBckFl+dm7MLX7CRWyA
2mf8Sp58tDVj7ZksYm8Gexsktc8xtdQbhgeVOmL6wAZXVwwfQlA0mmirdFFfrQhZ
mawECBu1ZqZDrnsELlVDur4SkVIRfw5bCvmue92rqVjn4VuMv732CIV+T8Jph8iw
+iD3JDhajXbBvoti+mqI1OhO0SpB3JAbOdN1Xs9WXpa1Ew3rNcgs0T5E3lZc2owP
6cMmmzb/MkE9LBNpVZfcQ7sMqy2VjkcEsq64wk4cczTvxYFVMsTnF3OLAoAbd48J
8D2pdV6uSPakQJYnGX99fomJk2V/6y6RK7eAGkoPCzaj0KjddFU9yrUkPk1p/kzc
LFnXaziZw+UiAatU8wy5gaejQcCC/may7RjRqmZF0eSu+NcF7jlyfu9SpcDVeMz8
mVvCwHSujBj/YpGjhS8BtLgQgTsQqStDnfMnvZ3NzImebSLDMY1jjQRnIPnxLNOY
yl3ltWO912o/rf/6RgS5gK8EpvG1/TFx9cXi7m1+JDuyoxEIdikHRXpYYleLFtvq
laHi0XdEx/LKzULd/Mk4tKwUGrHeZMv4hsbDhaw32VeP8QWDiu2I1rkaZpCbaE4s
tvRTwQXnPnVlNxq0fcVmDXVOiQlOh6x5/JEHw0QIY1eyV0vCsd1/Ki9Wflzvk8xZ
Fqnz2Bu8sUsOzdPMFiG5nQZvbT1nqozxizWQaoxuiqTOXuhafhWyi2e1jmfEWR9P
oBhG/qNRNwHBUk71BBDqhZ1Dpgr1XrMVL4WVmjcknGyJ/9gzPEdgr3OxjD0MAgBu
/nG7k84MmDBggQ//71j9bDYb6tV0X9Yx5KTBVXTgNb69UCjZeqlILOgKSKkl4qwv
+8ZuMD6tbX82a3GEIbc//itoTcXyK2YBx/T5ILxCIoxwPqBGgIJXLo+zRRzckucL
c8let5jVywyBcWAW8Qr7mbGZ6p7fGIuACloSIE414Az9aR4wQJ572v+C8N7sr7jx
utttTmaU1LX0sYq57d0CzBnna73ZYww8Dj6nOFcYPIuYxbe3aqbeVEEnomRbdXp2
BJc+SnOAxJFblH1wD39NJh1DoDOI6StKlgUXamjpHZ5ny/j6LBzn2U1Sp7PfgPqN
7F83U6QKSC7F1E8q9n2r0AfNowO7k5XXo9NVGllATwn/FCqK2P7JUAuGybKeTooz
QqYN0Jt8yLnAjAVUEYeXsrY5UwDQwC5JbdT6/dX6NEpSTOZIdAglHgPrAYIWquGK
DRr8zhkHmFZI5pf+5A0W41PmdywPVlbX1iB+7/WQISlLXwb9C1OQiATuVoYzemHR
bqQf9XISz54HaFVjKrex4U7/n6DzPIzJ01VD4Ay+Jq+DXwkhgEAUlqtW1PmXQRyR
Jk4FMA8Ya7ZYuMwplvcUaHVLQna5IsV390gsvKWgObptS2nJMSdbdBg9Et2HVTOb
nmtcGsptjfJg1kp5GsZHqiWe25Py61kcubZiQiCzLfU6EVg+dyDUeBOaKUMAnS+T
KvM3JNeGrmWdK+y725xRSacCjDzDUdggdiKT9zY3tz0fA/uIbF2423yyUbw/R7AU
ECvJ3EulodDYQLn6IU8Fp4Z5gecN5PTD9Bi7NEpdXpUKs9gMblxsPRppepu5+xhm
46vVOsQgPIoMu+8TEYuTB25fxC9IpX0+27l51o/bYH0NdAMqYha70adpESFivd7f
pkfpxDkkHhiOqW0dqR+BwsLOHZIYo8lMWN0tySRP09yShN06u1t1R8RvTNO9Tf+J
LLGHQkQXajQIaZ1BsjQof4h8LXrgOgEDQwXHWRc2zNZxGx3hd2KGGZ37TsK12Fyi
OBV60a9rRoxZD7qMjF7cKH9Oz2E5IDFsNF6/y8DRVoEWDXRPv5t95lehiRumsxDi
p3Si+DtIkYvvSjoeuHv82oB/pR0RCld7LidnQTvWmMnF8Axf2krF8VTdpjMytuMI
Qgfat+QG6n6J+G1vuzTsYa2u4xX7HI2fD7x27xrwzZyPQdjq6/Fiqcuu7cHSrQ8F
WYxtH+OD0A4EgR1eULlhFdZXSF4/Y6rfmpuL3N4mMOZWmtAkx0ixpf3RuMb4N7o8
/3x28d7hwxLGYUNYJkxeXhMROQtYKIFchEKnhApENC8QE4wOC0Hv84GDP/AHBaeU
x04Lu6OmEN3vIfNQnGrv0hsOja3Hw6AmtcmsRjNNj5LjuEZ1MI91WBjTrnf+TQKl
P7B5kYH5633L8Xx1+yjF7EMh+btAbn+fAQ8FWE9jDCkABJe8Hvmanc9LMbtObXY8
c0hkXKkXSg9m9JHG9bNGN0TRP1RPsN512qTipaYIyMyxeS43HEb5/P5aKvtRpYpp
Q6sEAGAJo7x7XGo5HmRHeD8A0xOH811CEIgIGJ71yuehWkdtAPrFdQy+kixgYhCD
RdcLNc9A7/DmBD2D3tPIczUdBe2Kt+XaNs6vo4NhrFH0+obp+sM/skDM1JuGXMZp
SSPKfjuPhNl8lEVnY4I/cY/LZ+Srex2AJQABhgF0pAqcbpgs00IS4hjjX4HTeSDv
jWNsDAUpes0RVWlie9zR7tH+LlPoQbp6aucQgPGM6DeU6gZdlHOUBB83ajeyRUh6
awBMhIYgeBKgD0uKpowaKaaDYZtCc9N2NQ1uklskJltzyzOAkiyROAqD/xyPXSse
/p4r8zPrsYAiEYE4QLt5LTxUAHLyH+/oIC5XkVcJx6ZmgasVENSwMpqi+q0MaAOe
xyGSwA4xQIqblYYZpEdNADqM/sQnHwpoJ91SexqDtAcBV5i0VqQBbN2QspiBImpD
NfEVKzUI29sSu9zAW22mrMr7xFFXCLfB39Bss871qaVZecR1e5VwzgVEUJpRifsX
W6BO8fkkEvHsY9JRyvW+Zc+MKGJPLiKR4AD35EHzvCpHaIVD7LwvjHRU2J5Ne6vR
B1wqx6EoeaX1BSKDNYHRKY3GYlRVXfjNBaPxAPl0Eb2yCsiXi3fglgpV7JCWeqKs
+mV5e4i/NH6uzMbWbfZezCCaLSrxsJyMzmyPBiQiCC1cE7x+CCwxvTco4mL7Vge7
i+/l7R2nFao7+zth9STn7Bod0StFCXNzbovJFB387ObpBDwdCqOXxD7M/W8r46/4
RsgKpJkAJLMtQcDbdfvP2J98avHdPuc1SUU7NSGvDmSfgv28vex/d0lsUY7Qh7EF
f2tokBjfHE1alEqilq6sHukwqA5qFZpLg/+ag2Z2WJEp3CqxVE6YXpq5TszNVBM9
8RNUTXjdJJdbOzFrMyRfqHL/O8CxSoGm7qhdA/lyUEJ9cYFWVLQ0jLHzpDE6r/lG
p33TcICsLAgH9My2+iG/T0ggwy2jOdn8bsY0cRfhs7XgpyeXx4iBThq3h55EFPNR
j4VazFr5ebUVKY0gGXBuMGoSHfcFlYuAmDhuwOfhOpRWheRfQLZMHtJ0RMPZjEl7
jiz6rCX6q75JOqASilA8/HwHcA8k2iAbT1N6QwL4k9b7V0jl0+7RF9rhXua/G88c
SPIEous9dzja0qXsN9sGLoNTq/HdClCtT9I5iW6fLSj0Ztb64PDNggre/8DhKq1E
HqizEPpHPCm3ov9PlurbDp+dwGdOqQ5KJQJMnqbP69zed6UbKSlaUV/istsumeoM
oKr9/Zt4x5PjBbJJVuu4coVSNyhkf+4VqAdUvs571gOBgeDFJsYdMGL26o+BQn40
jw3oSJ51q9l0ctU+fLS3ngUOyRy7/eyBgQqcbY6OcLR7n0AHCYCK3ueixpGqZ7Zx
GvJ5l8Vv4m0s7SbxM6KvWtTfU7zODr24lrWYC0y4ZXhAuOdHUoyn1amGnmiKci1k
3X1FEHqTdlSg6Al+iDYIEHV1U05zr1jcsex4jJByP1gpl5NFNx2UsuvNUhErpYOG
qNVpBQXZwuKxEB8sYcGRSFiBWLJIMf96njX+vWNZVyTVrH98Uq0Rv3VDrglRI3MR
Hg5loRVWnTgBeG7RitiK1wkX+Itwtbh9ZN8PjI9d777A2uYwnFlf0uoNOVeurKED
cBy+t2e0F1QDdYcxrJjsRVTQi2xAz8znddvAgiQwBtNA9IQo61K2UqQN2r/pglmQ
mypemklY7yiS2pcHPRfzlZdoLqvuof9Sg30n6DAId5U2sMF2IIiaA2IU/1Kn2R4m
CkoQP6qDpRPqn25hq87vELBPOnKXnRIvB3E4Pm3pMH66OzCS+rhvQPBcwG/p+Eo0
EnwLStxuphheRzSg1j1b1nd9ivjOMtEncHxiJMI96jRNXr5ZB5LBCcIt3e9srZbE
46bpXMSX1ypNFnTv6Cb+z9kAvXXk3sxK2QTJ33idA4eLzk6qMgnBN6m0+1vzDWkf
9xQ6D2EcZB7khECDAVuPc6JbQdBmNUu/rU7DcRPJp7lHcGrXj34b46gDQhRo3+cQ
pFiTG7wkT/NQ9oty3iJ+5N0pAbwJnSTjLgmFcFeQZ8ltrvxcRvb2rNwK7bDULyPr
DpPCk+m0Pd7OKHIGWCzrh/EduMFifznBxS6QENauWvrM/NN8LRS1wzOtbgW0cIZt
1hYkRcuRQPavh4Irq7EeDLEAcUioqMb1MibqMlZ+/+0/bj7z6OveFJ63Lwt7JL+u
PNj7V7Bz8P/ul9BGTUmGxf1U4QP+bM7mMJPAEUbYf+fHKXwc+yXcnXaWwtRYzUN9
zFhL+0jnGxSdcKaK5pu+JPJfw5UEfahcujPDmh6ISU//amY7FbyBUSILv7Kegr7q
S7lHCxJVtRSXdiQTwptz5UFFVXBFLodStlefKEpIEn0uiJO9ihiyH5l5DJOEx0dU
3OgQFMulKmeEWgbTLPm1vtTf/x5rM2nu8QjhTVz1/B/crnz9ilj3WN8jh62Y9VQJ
NtfL/PgIKP38Ul15p7aKPsl4YxNds05q0fMwW+3EmpsNVb3+G24EIBPC6bsQ5NeR
apSN3mLvDXOohE/vc1YXUgUL3ckdhRZbDW3j836coTpG+uZCmeEO2DRs8l9WBVmj
8xmqP9J3Vrq/BkT+gH1kCDNADJjSzzFz02wI9ok2GBaCMkbkJtEn0MFfXqQSjP1y
ggcaAr9L27gzMix1J0/4ZgNMl8IeZ2Z1KxwwMp8VI24Gtkm6lxGFtLsm1R3VOhL9
/JVdFG/upkC/pKyZpWt7/6pGtRtVscuOx8Hser8KEw4lRasjHd+LlzA53cjBhtVF
b0Xw1duZiuIU0gNjpFVgAEQ/xr5lv4+JKK1CN9KavyqQmYYzHBDvKa13Lj6JVetL
60gQuYTkPwvyjng8tdBVNKhy866YSoRYncJ5T60XuOkvTl31pgSig08bC+evKNt5
y0KAPmTvTlvy6g+G8v2yJ4LCkprKeINs8T6Wnpl/g7j/VqaMsSGtcWIPhdQnYZ+2
z3QNkZ8RwZgG9C9azCrGb1MiX+DeQqI+iVmQIs8RcE3Pk2vfWIfhIsWR/4a1z2Na
aVQt3vglxIxUvSdgkjlRSxLLMfwxPj9DCt8nCjcko/p92E9fcar6qxGmdfsWAVrq
R9gokLkXXXtjcsZO9y+t08q9wpxw1D4VUzUZu/2MOaWfSpreiIdUKfTPC/Y+xVjj
Wc0hZ/I3mKWvYL0uNcyRZ3Yz+KBVvi8E9qJSFpzzwR4vJHUEKKRwQgbkUCz52uO4
zBeh/vIKE70lmv1Uja8sBuyopcflpwTer+EQisu2w/UhaNhTEF3PbXXSmvtIc2Jq
43zHgvJSZpthWcPIOOPpzRk8AzeAiGk3pCH5N8lXie8tjVkkMJErsGaYAYtpPU/O
KFdukeHUjIlA3PT3klVukHzXAmEdV4MK2bPlo1hAaysIWywpWa7JZD228If5Lcc2
65Rgc+be1sc8CEeRHZH1D/1aafXAPxH5nfPIJS5+kS8WMByCrbeL5Kw0XhTTVxXM
a1nCl0h1fuz46tlE+7SnuGTtGEfthcc/1nEhSCUvAlvGNocXo5Vx0bWbdA1YleV5
lme7tqVDqnjgwMRtfLvaR6/gsD3j6QXXEIcnlixcSm8XqxQLD9mj8lu+0BnLTKP0
ECeOaMchryBaLyqoeRcmI1EpJfscwgKcnkZarb9Qu8Lmerz9MAC/pnAl+oS0iCfL
65ltZGL44PemIUJ2bI5gCMxI4GLXU8O+zfEnHmh7P1u5wg5BnI5sfForPsrKW/Dc
K4FL76Iamk2MH2+lOjENgVQpLd1CNEgxTk7KKoUb1rF4M1KDbkats/qrcTq9R8H2
W0evw3tLKERJzvH58sbNUaT5gf6Qc5IRBTeGw701JuO2YUi90BGaCtCDcutjiynH
i8YWfyzW9EhLNfSffjUWToPeYS1JbulHqlD+vhLCsRpzxSyz5JP83RwfmdAfbXw3
kLCIyjw1K6T/HYf4s/C0yG0yL6Ii9D3LrCcChlvD59v0m3hkcNB8nd1fZxypID5C
S7+zstwsb5JYnTQbsLp9Cw==
`pragma protect end_protected
