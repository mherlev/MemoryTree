// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
D4nIpqI7m3miwZeGcIpyz0liIymZfRxLXG2nCMOxEb0XvGTiaWIzk8hkI141/eGF
dQq5ctTx9Iq7cbezG5ZaQUCSD5H5hfHBOSwTJNySjA2VWQRZRAQ2vCcLt6Grf+sV
/wY20gxBGbh2IteuPExcXEHseKZ8ToQCTY079njKooWomErKZdye+Q==
//pragma protect end_key_block
//pragma protect digest_block
xBd1Sl8Q86AnWkRhmP3p/RBvlcw=
//pragma protect end_digest_block
//pragma protect data_block
x7hlvjQfrp0tY9rS9Dizh0MH9VfnfeSkb8mirPylgaTzGu3kHYJ3B+ykFddx/kS8
u0cL7RHfaK9UYolQEgsRYASYjXQ6KDPHmzUw5ktXk9y72xMf/bLmACw+zOUHasRe
CMjuX3Ex0eJj/xSgIw8yFzgLM4bk2liB4wW2co6vUF9ddZxeK/M8H9Ywt70Ug+Ta
P9pTN9JxdBgKRxpvPtuXy/bJ0GwoO9renkIib4AE49Ge0why85zEHhg0jS6F6gWN
6pGXyWN5AJdECKUn7X5Ao4NqqPZd7YJLSVTBxdBWjhD0H/aR1s2drFvrCEhZ6FAg
RWt21cbthap80N3KJXx4ZCLjG2ImLgnpPzjBz/g14Bsia0nwyThJhnT+u9GjQlN/
e0gGHFQ46gwRBDvFilzQT4WL7X1cm6YeVfITSW7XJYLML35lQbLrLW/1W3Tz8UdB
S+vBaudKpGv1qYxzKN+9+umnhd+3XPb2fZHfGGoHm38wSPNOApgIt7RaJFzTKhRL
e51lfYLwo72QygGT2nKQh/WoC+ERm9iTn5AL4eAxnW5MJTPAgL2pBBnQZ2amDrFk
cDkyAZYa1+woQNvqb6DoiGkb96oEVSUqDD8TzH+60R9ftbgmWQ9SJiL8lSOmKep/
clgr7uULa4GshM/BiRNDScbj+sBdONXbcPdlwx0W5igC23FYtYyIYiIBfIK+FWdz
/zDo2CRY2MjdcDRbTdT83dZ8Gn/EDPuHUCz7coN8nhoQ+Yk9R0yzl4PUitAbm6JM
iq82zLnBGqzpCzzP1R8ejvPMxNxwIzU1PHYn5d5KzkA6usisFrXlKkWNNr0DOjm5
I/LeSBkgFWJlnOrUTdgOCYC551RbJYrX+zJeJpoQQXQR+Okgl1BePgtM53sR3YsA
qAJwcTHmXUw2kbSCm4dvemnv4ej4J+K5G2dGnaS+cAjtE/DXs41jRTze4cgUb3IO
x8iljFWG1GHJQzb5V4tlibkteSCfnibnEIcC/AgORdkS7ndyJEQ4KKnGuZMeoGQ/
x3tiwkWtUwgTYRBzbQDUJB4POHuuv7Hs4hXWs07H8LRpekusanwpuDhGGSV2Ldpg
bpUVXcetisOvuwETHejBYk/5GjVYvRR3FedcpSoxzo3zb39F+tZkBJbanXQAZGDy
J2jbHVzmQUzoDOF194yEgjhcVNRnquFU+FlRB4SdozoeyJAS9JwRxchjduMbNLlo
nmfRa9v3iTjbFIF14yJ1YCidaHhyNtqYqIIvw/kRkryaY7Sooa7wqzCAzOee8ubK
K5G5p4Tit7WG0eqjFneyArjNOJQ6B3MeqUjYtK0Yn6G8SJxviWjpJ4ogzxxsgmf4
6DfLkA0VLS6Ld3nNWRFqnmOsZENpaA5RhgHerTXdWz15l4BHj0XP0vK4VbbJOLyc
400lDMKQpAMhwBNKMS5/KRcgDpm/6B3dXkzJSP0E7S8CxiAIqT5O2t953N5osaYt
1AwqZbAN2TSfx0atvwzxH0RZp8Ey0tV/NOznyaoIBq+q/QM1rHnO6iCpjOAzzt19
KiGW33j/dOqHEpY7IPz2THGlSCEWuoBqsIY8jDUE2HA7Lq9l0IB77NJH7z99Iamf
ndmQM7LhWUTVepY1h5sL7PCnhcOjJQxtaOJYK2LSZdih+3JnLNldt9pyaB/4ngSO
pDMaYZa8Qn9xwtWR9QfsoXfsxwNRr3ju1K3/XNkeMzgxsfZjLxTntg6zBECtbFVI
u2eKtZ1gxqf2CaY7Ru9t027R4vkDPJRRRVC6zDORuxY/M3Iy1tqsPGfrCsI1P0AA
Y2/YXEaSyrzwABiVTdFY36ZW0+gT5yQ/S2pJ0OBgnYaB9ZYkI54oacyKufUOJjfK
u5ZWOdy37+XTJJUlFSEZbisZOASzMpX0EqNYl/9rxPsBHp9qmrSwZPozLAV7vZv7
C7E5vjybbFxz2VocBkFlLOgWNpuXNfwYbVrSFPTBL7u0OJ2r/t3nZYlOERkBOSye
JvuHSNGB71KpeZVoSvXBek3/FNVpyBL1ds/4rUrC0mPhyjqKcPbCu61MFIhlTQEE
hSsTb4uKKgfveivNRlEuXPjdUMIy7KJtkVoKCBWK1sJVKdL6cgYjRDakpABtxCc7
S/2dQqi524Y1PTYjW2YLK4ecFtRR+K3KSDgRXu6SQ7PLLli3lv9cLBZYNLDKhxk7
Fvo38ga4m77z4x/yY58AEx8FAijqWm6T50BPxW3pVLpE4mXyEs8yjSwt6dkTEd1Y
mLy1ogS8OUb3Dg7BbOs9TgVdGRYO8wwgZavuzQrvPTzFru1vSb0461xV6qkk7Hn/
oKm77CNSHhofa0z9p/vuoM/cvDI9Pl7eqbnkcPHLHNKPfHDyzSRGDooGb/ShR3xp
Giw6TSGHxRImMZEmmd/jKENNFCW0OA78SJo1n4rmDn0Uzt7TMs0QdgmVe4IK9nXO
nc9wOSknosOIPhrZ/iq9vnaqATj2b4x2T4jdkHYOJZPofO7K5jyB6cKEKjAqpfhQ
leotR3q/jDY/C9GiIQK/pn3toqPSQ/rwsSxNdmHyOKhyTmyK2zen6yZs//OjBq4q
z0mXsii8YfzW91/FE1Hia4ZvruXp5bmc8SHGaJG9FmAbZlYrM2rMt8alIfGLvg68
KZbsbQzUmoyO8coU3SdfbMwhQFhtF1gVl26OB6NLkhLAh7fQSHpEJGt3jiwqP5ab
JGDSObl+76JGusVw9J7gTIBGY7vQajNAxxoD9ojz6aYUMmQtzJDeapSseUj3JcTM
m2NPdI1Cc2qhItMeLz4T5YdtBtqbgXuGZ2r3mcvfQtWExKb8zAHPPS3jWyJyW7DW
esIHQRgOvjD1G6AczPLXGef/aSTZBA5gY+hgte1Rle54X4C97+g4r1isdarmLNLt
tBPortHhvsbQcZ7RIkiGWgH1Z3a9QAHpBq4JMVgP2uGaxXRdd0Vj/mpJojcrW0Vv
cGeRwtqEn3oIiZLE0pbwqBia+GcZBd8QgJOQAC6cxrWmgbvP5XmOevYQkpryeGZ5
f7dOnvRbrlXr1XuALDHitxVp/5uCVP0HUrw3x/SBlsTV1fBWjERr6i0RbU2VYXfh
mMgloPTxiYOyPbZblvvs3i4ggFAlfXKEA/SxgdIFr00lbrrWMMbyhJ6at6hZxspL
GeeGWVp4gCRd65Gzv2NjtF119O86P10LJaEl7jcQ5Le+4E/K6JPJSIUiNOVpa6RC
KELh+oJDSCpAbwYUQmNAQzBGRB1XkS3bG9sYkimjm9j4vEWuc3JHj9X6YzY4Kyw5
WpFP6XsGQ/XVKXgJ1nzxYFq3To9pjZliijAzTECEjSLzd4h9D0hdJ/uhDWcNXaL5
CjX6jCs/hb7D0m16d2x534slKlZGO6S9uN97O8oropqhI4G02ES2cxbpoCIW2vw/
ULNKLrUYbz3UC8j/Os8Do58bh6lfig6bVHtBB6Aaol8Yk//z6JAzmyfJqujDoaFE
G+jTydUhdEB6pEyJ3KQi9ZNlvbO/vDBmqQiKbgmn5OLWUu6cq24rcOzDu21IEGZw
1bIjTWJoqc0JeBqHG0tr0ZXTBjThjAS91lFb0ticuX99u1OWoim1xpIEt+zsoD1y
0vxhj3PFySsT72t9iiupPIvVnY0JOURdF7jxuCLSZZ57uxAbbJuLzuTTRjAb9bLP
j4sk37JfxRJmoWzX1AsIopN/lv6SLR9SCaEYJKsw5WsGLtHu2quUbNb23gK0H7wQ
FlXkVPCB9uOLtz2koWydI3XHtWcOMsuWdXT28BB4TMXsYLP2Kgq6Kg68jzAPTZxg
DLNfGeHVK/laZ8Xjoh8SzgMNUkTypA75xbNsIUu1h4+Xtw3DI0ObwXj6fJenuevL
eOXqP/USk1d5unwgAUsYbEckKV6goSROgZUPltPd3dIytJhf5WcvH9guG/8Cb5iJ
yqmRia46Fh1UrSogA2kH1Fh63tQ+ChpvMFirBzkLf6djGOGMeinQCUDxG+RFTLTB
wqOfjzU4CIUbcqxTDpXAqcYLcUt4XGk/MF/iqsTGijzHBfEXAckdC0UElM16/K8U
+Rie8SO4+UI92hb/I30MtYPp6TPBkzOwYU6u2jHf19V04Fnmi37Bu76yJbstY5dU
+O2c539i5FADGbMMbw8grKF6anahu4yIo6LQ3IIdUibszLl9UQMlmnY4S6ZPxeNA
H2/RD5tMu3ERKw38N+7bJCwoTphbS2F37h9t3dO2olWXBj8nozJ/cHghZi9yWewX
tU3y3VAWwjx5zo50gaE+t6wVaiGMbPoyw23qVM3ZlnixsocNUX56azCDhB6a5aFu
3Lq3W+pXfKwnfoyWHooGTMiI+D94fRZHlhmr8G3Vk3jlgdzCZkR8tt0r3tRGZpPs
B+F98OondhIGATtfF91VbZVaFKBmn01U2R3+oMGKYKhDuSTZVTmMRxrnrDMfumm0
zOJyc3Nnjzg03lVFH7pmWpXUP9V1SYJfLZUE3j9ZjH+zNbyuZYHsnj20e3/IHN5z
krb/Tb+M//KJ04aIGYvcUFzNdnwSf2YblysZCOkAT71EjU4ZtAlk7AdhXBEtsasV
irlni9M4ZmK5w64FlQS/UU1E5DBWJPp+pnaLUIwZjJLrxtDkFfJny8SrDYwEmE8t
4aey/PF+Q+eLJUn6118V8jjtQ1+c0rWyrmk9R2wLQFcPS3XvrdwWYpJQ0wXbL6GM
FGFTUycYgFfVQSXZkiROa0+VVIaB2NuEEfHokk/38AdTe0QoA6Nca6e89PO/WWxa
3ZglTlUN3EzcnaDFdNYh8aonEaynP7ia7kIlE46pIntZ+3ko+OWCASA9fFsUCvD5
WrJZ8g46xM4PNhW2RHzA+Z7BNY+F/J07fJYvseUFfWXzjzU+o0k8NJAwjjAf/HN/
77VDA+KwAsqHv+ZXRzmtlfIc1PtjaCpmMFDDcchTKEDT9m54YPAj/6ZrNiYWPVwY
T3BO6xEAeDE44E8rOKwgWkTeIUc7pF5M5UjDqWerHoPTFlk1XUpKmVYfBZU4Xp2D
HzlkFNXM1FS6D8RBBHAm/LL25Sf+FS7ItT/9ghknRD/zzhjDeLTz6SakcMW3cDSy
lfrKo0ZlIob+Dt0ezyOsouj7x+3nuSYJ9rMw1nmDktc58JpaWmm2LuZKHBOU70E/
9ksjRH8qr4FWXP0jywcamyJVwrP2W65siljwu61uYXZmQ8R10d0zAJ8qfSjvmEZT
E6R36o+KhyXIYbLPelWATh12soIZtqcYMGYez+yBB7BfOp0Z7LkjfTXExblDsTZq
7wonVDBjKvcS4tGP8Rp4Etn5oiMXYd2kwvfcoX0rYQj3+i5ZqGY8QbsvwW9l4Iy0
8WMMqCWTNjd2ryj2Q3vhk1OZlbl/ZSRW17IMBp+DO0JeNtkE9EUGtywLS3me/nGl
H/DTrpV2DBuZtgRf9J6Xt8NE1e8qOdn3hpH5up8nFeZn3XOGOMmhB66Z5NUMvmzH
Vr5/IJJWeRmiuC1P9aeCB9swHPZVF2fXda3I+T9MA5rfwCFl6xgy3gN2BPVdUGo+
kN7Z+Ex7UPc3qYiTF/zKM5NOPS2MN10GwF3HxIEzkuqNXq7Iw4ijttY1Z5hMbvTs
G4ORyw/E2RyiE//QJ2DO2bDzAW9xHwcg4eMIKHXnA5IbDJTeCEzbBOkradJSPagF
+5rCULhp5StisCsAPc9XNtmPyY28DA6dC3zvxRS94zfn81rw20W7+0WskF32q1+2
ObXoNa3c/7IlhgH2SBi1j7iAkuyiXQayf1G+lX985Pp3LKVnLuvkHA7wVckC3cwu
X8bqKu+4oRTljYAp2SjMOHrpqw1hgnjYqtKl1o4Jo+XZPgL+kwumHRLPq7QbELeT
ClDLYQgHGoH8j5hWYUSHc19qH9Nje/gAlq8WecmyFCZmBxW8vpsKDaOTcscu0BIb
R4SqFVLEIZA3E0f4G1BIkJIqmacWvkql3r/FgLa245ONq6hn3KbinkF5Q+2ToPEY
rfenYIAZ/kJnaB2saz4uE3Cwc+gcOpmlJQd5uxpWNzfQ2VjYIiYij+YC6VzgJ3EP
48SLJlBFcz8AOf0dtZsyO1z9iSyVMvcrQ9R8gCo29JvGR2VHlDczMneN1kGEysvZ
4R+kJaHaSVVfr8WLNPBfxXjU4Xi4RFU2cgXnL+oPEardQ0I8/sTedJQaZm8f5gEv
iDhIsY60oofjFwWGD1oHiAuWaNfwD+KWdVfmPfpTnBeB4rKNnBky2XQXGzSw5VuH
ehFPNWF5SOby3pxkCXgsjIcmE1k5qOSKO6U6/VqFVXhXtF5Q8ZWKLVtd/uZOdzs+
y5VkuIgfGS5UINZlSaAu1W81GxLJ9erBu1SWaWyu/jfBTs/urwQxhzJO7EjEVL0q
cBfsKdJ2iiuXt2r0z8CNYlJ8EoivW+LF5T2ehET7w9T7w8u+3G6mW9waljYaY3l2
kkc8MaHyHqRE63LXwWZx/xWiydqQ7/GJHgkxg4OlQlAVbYGjSWdnmJJbXyeDESeZ
txYh+Z12Y3UhzlPB8B5VGB926rVe3MHaincPYry1L7+GhkuFRIJdoqq6gqappcPE
qO2s24ZbaNWrALK7g0WwX2pMAwm63A3ulcIBYYjuk61PMxmKfoj5Zef1I3za8Hmd
gaHXoUJSAO9Dv7o8BrO1HIRQs/RXx2AKSVv/a1QkU4Q5qPzJSpl561noUf0i9eWP
t1tZTdXx27X4w+nXxJ7RYqqpLhG6N3LNLtAkye4tMZiAdKlJVH2Ui+RDvzcl6M9v
+2hl0a4SfhKesyX2QYiDBgswoCNoYxDj2zfXQSNJGBF8bAyzeksjaLI5tbSwA+UV
QOcVKlxEiHurtkCHVWvDd04oXSFdGkb4nC148uNnd3yzMFWC1JQ0vL9dPUp/OA8B
B1aQX/UN1l+Ltvt+BpRbgZkZaRGZ42xEWNC+a/mKm0ZQHAMkU8Th07yIAwrZEJhI
5Av7pycxRZJeL4TIfyfQ5atmY86w3ZFGMkicoKwlMr9ZmtkRhBw/PLB4stDJ6Wtq
1xx6wEXzJJh4eoL/WklRNAJiBZcnZz/JQ99D6fjrBpKE0bRoZh7jKoiuRiMMySHu
1CE/guuHgEltRn7KBSDVufZzO36BVlUzbaQ9KgkwW9kl2TuWbPVxgYVKy7MsXS4D
pgIhgCIDpE9wNKPC5F4IokGXIJ56ZKdX3W3EbUn9k1xcbSN+K5YzALe9uzKnUoo1
/XKVcW11nCvF+0RA6/6tDzqtUnPpyoyo8ZwWOVCOi30OY1Hq5fD+9WqLXz2Z5sb5
0dSxpmUHO9NyerEI2loxQi+PfjQqx44B+HvDHw253EuIblyZvgnjNGmWxKaOKZql
vguBFyowBgR6db/Xn7dUH+MwL5ew78OGGBOLj+Q28x8s8qVnwCQ+Bl1ZsclTdG4v
g5Ufb4GNHxzAvQVXpwj0czh0jTRs5L8fk0EDDWjJJ6N6eWnmb9suO24eM/pIwQl7
VoCthXSsGoyfq2/H95Gg0wV34jk/BQkcVmF+ALrE3lt2IjZ0YhYsPT5Dv359m+Dn
sR2efi+P5vsgWw5gIqJ5r7Lv4oO8nP9djOi7MY1SpEnharZvC7Bx01VqDk/0DZYF
CX7QZ4lJhab2JyjF/pApMy/55fdLwfGVwDSR89eckHLCzogzRw9EisFsxDSgVxyg
2arxGY3lmHZvpG8VZ9H+0Yu7nyIZTS9ztcgzOtF6YjhgVnhq4x3xquUQvx0RsJnS
uHO06AKcz3FroHs3aCqOzezqBSaf7ae/Mg0t/RKGhhJmWxVXVUgZgHZsc4IDkR1p
2dJKMtZ8s23HhfLZ1fJy8D9yfKi/wUU6SI0phksmtICXG3pTzxWr2lsHq7k51UpV
wGqRfBkYqqd1tiseekwq0y8RAhoJPQkMpQytA65tXbj1VkXghrEw7s/1B8RQ8aRT
Mo0rtAq9scWCDYJPyHKs0ikP2DRI0pWj15TKQ9UPkf1loyigE3ochT4yQuYM9voZ
ZkdjZxnibkUQ98Hm9dTYXn/gnoQhDLg9ha6AP39QUd29uXZbvt20+AmjhI+P65h3
hs3CLPB7CiUrXdNoHj4TJDHRvVeP08RvufLU6eySr5n+vZobtZ6wYRpwxydrh5HP
UDNQm9sGbONPERKLLSLXBdDzTctVLJI303uW65Nu2HOv0ORKfGoZqf+JV1E5wVqi
JfC8Sc873j63eybhTSoijPgnX/l/I//ciYisOgwS01hDIuu0AEye5Qg7dGr8wdPR
n54yawaLrvdA+yossiJTBnhBtyMidvUUnS315e/y71xrzKU/V7IovCz1kXuO6C/X
rIdrtNMoXGfhNafA873LY9/8tz1if0RcNhM2BfnSS1ZBPvuKbfITRXxtSf2XRgwk
Pk7IP+CRLBOT4iDKJ0tV0vINgishX8B0zV443eQ72FU/dDmnBFwwDycHZDTZJWsN
uHcRYdLBhyHmDtKNcFQ4BwwW8AMLfzqgEs14yVyWzzBvB554E6gLUldICuHT386u
BceQXnYdMU8Hbc4HIgMfsBj1XSM27NxhkxhqK3HcjyfSXphWNO9ZhJcvzIkoyGkj
/xc3BLvyKq1SqtKhrWFIrM9yiKwyA/CFE/1n+PJbztZeMjJdms4fiFw29CxipwUd
z4CcGApxo+6O3ALDjudrJDnOrsaMwliPSVlzsja7cnGmP6JtUXtdn/sM+Kce9ExH
Rw5S/UraW4AHbaY9ev1VJkjOvHtkL2rLpG+P/ZYFNXPw2JA8XQJqUaEHUR0K+WzA
cTOWMidHSx8uXSl1YV9n1aRBUEQDPf/Sl5r/dCnCBCBUlzU0WBM0P9Fr9zZCmByo
3Z5njosjPS9CZBmuuotNtiO82nqcS3c72Au7ZFqr7m8rzqDVDGh7gIwamqBrwsAc
ptZkZclspeb20b/aZgXVGVLZDrRCep3I9HSpUfXxonhi2zOs/tIsdhPldLlRMquQ
d8g8Ql5BJKYEFomUPC4cZy/ewTVdJ3jCDbMs7m/js7Y61S0jFoMJsCepfCTHBVIb
3CULrqdblox5SSooLX4zViyzwILDCgkPsf/RpOeBMsriOdMK/aYjMwBh+MMVXcUm
9nT+CFup+wGRlA6idGK8HbyeBdFnIoH8XXfdoIHtSLpvcCGPZ/RnIshqJz7BYukD
GuOvVAIXmMR4LNMaaFlPZ03eP+T4sceTd4W/sBmBbj/3tGoBve1QIWwa5iZv1dSq
mf6m0eNxfabvJPb1f8+ojOraD94MgerHgrODLBZmLr+gdaUlYBl5OGWbZltne7y7
dogxVv4bMGBvBLYVYOGZ5n7f2hjgEAagyBi74PZZrl1V/dGwnNY+ocyFEWw+jem5
LGtVgejH7p65iZV0EOpk0z+AhdiOp4FgtGgpPhKYUDqbArYjE/UvErwpi/vOVtBe
EC95b1UhVxK8h4x9pHdGuYSHNqYEXBaWJxPrGn7Gwb82sTFbpXTJOW+Xq+gec48N
01lWMdzpFi28k+oMKCKCUAkVyzko4a6n+d3PDzPUlmAQThckOn3qakYwYl0P8Ej+
QZEXm2bcMixW4Y4rtUOe8K1H+0B5kRfw6C9KYQ4kJ4JPCFSO8yFGATuACiZQ0tIs
3y3ji7RKfnOBr3C9pkI8gwjMMFafVRfEiHmcznh/qSTKoHWdnE+ytVpcJcZIUi8m
R7gsQsxx5IgtqHtF9llRHEoiaGQclxMG8rmOy+k8CsFv3dN6gKTCOpPxXTlkC0wA
YBlAsvXYsOEu1AHvzTehI7XJABDvEQ8S4R9o//GDT02HjzXU0ZtnIlmnJzcT7707
zGdaPcQsOn846s0TR7RtaeEBDMmFRA7/m5ZCDIu6FKZJmSnt3KrM6AB66YVy9nGZ
PV/G/Il0jphGmno11KQw3q389fffIQXu2tHkITLAGaCmpAPCJ7KDQybqlmLzogRp
CZlG5z8x6XO1FqBo38IlS5LK4ss5fFmRVbt7Hy4Zq3oX9ZlsMtsiLTR11M/gP/dx
kNSJoN6Qr7tDLTA6FBBhxxPx00f+nSP0Dgk5MbEIGVXsQ5Ezjz8eq2kzCykDqC5J
bGiGcN7LYYMlaEQcXGw7ad+WXCDZZuUB80yMeGcGq0YfsagR8I3n3ezvDqH2u78R
dxWyfKA71I7AtClMrN+ZUpG7pmK049CNo0SOo2gfdEnFUKj/nR3nHm15agZmKHr1
Gy9iPCBon2dqt0HkkdZ4NLCbQt4NmVUPKJ207dIIehTFXF3ofCBMhfurATMewnXI
4s8K1VTHtUNVXTKBBP4Nay9BxiqpoWazdSlvalKVOBOV/j1lC4kVrwmW6davxnO4
ThTzX6owikOnIcKGDeUyPNwvPGuW4EiFV1BIc47iZqBvjahRVtXYFAa1YpmVmlRl
SAsG1mDRB+Dr7dGyl0CXp/Rni9vwUiRcU6S7SlRzTtjqcweCmvdstGJrdaErkq0d
AKQgqemtwodRmoubxK0Rl7t8Pg8VpTn5XV3ht6vLe8DjlavHDv2yPR35nkQyXci1
QpIcsg1ESwauZexk2vsgxN5ndS3IDyPkd/19qEmTEU09mOSG7WzrlpWqV+NIP7K5
SNAWVEtaaHIQ5G2rV9UM5APRAuuQQ4eErMipyy5SYMJEI+CAi6lmV3yAxs15P359
qJBWtf9IweioS4J37F3JmOXwah+qczo7OHQJOLoCMij4Sx65mUqk3RXr9S6kERCm
B4buIgzEPdMFaf6Uu5Icvl6oDtGkaW3bdPW9T2Xn9E3zp5zusc9ploObXw8fLoxN
XRqVRIFeTrsOKczOX31qYjkBDpTAF9XYvCgCi+GNpz6y1/v/dk/rOmoO2jHlmOqP
C6DMe2FeicItvQci1qAxaZ9f8VsCpGyIfDiPIFCrKHjFqLykJTLUw9O0yikNjpic
Ho91FZhzm33Jo4RnJLCbKwwi05/BXa2GkoFz4JEAZxJr/1tHQPdrg/zYXWBaRh+P
JXmYzEXF1v0HtyOGIkj5qKcx6eLCZgE/FDJSCvj5+u0O6Ii5bctFFk6xoHgh7UeM
iJlUM0Nl5GJXm64nIuLo/rkmZHKYrimgFEw7n+ua2Om82uDD3ml93XVjr6HcJUFp
kyxAOKRnrjSCt+0K34vpFmWbdkW+iQqSAhe4IYKrsOQ8gI1872bTn02ic9wqDzl/
wsba+/YlDY76LAxFDNp4Dmdohd390Qj/9w7k9vmIT7YC+U89KSKbk6+/xCqLITP8
mejIGEzvnB/iKM+gzM6+Ve6XITjabGE2ODOBnXHNcnqPYSXzB5TP8PrfMrr5AHYW
Q2DHmSJmc5/NljcnaGAbyDEiCIayDAs4R9RT6tWqaqWhYVwuekBFWIzdD8XjbY7E
OGPTKwWuqCq7ZoJ8SYPj3Meh7EL3AmIDfxkXfnxaLoAZXY+a3G9NNcrxBETDbYfg
ZM51OJmfYKL1T7vE+wOGNEDdo2CrQmm/AhrPpHcey0/VfsTZcSv3CutAamk/bQ5F
0kGnsho1mfmMQb2WXb4/V2CBAVfztpX6bz77uiyEViaORres2aaz1xL7WnMMplnK
8IyRMLW/Ze3Ioi6jDir+u1sXzIN5G5mO8PWiTkVVETH9plOhWgxfFLfglgxcdo7Q
cn8+qO87iV8Cv63n2v8FuTPcazljKKusms/i0hWuGchhIrmeuBt1gCp5Y0jSSda3
EeEipCbdZKZsYbeuftSabcS1kPnNU1GOLjZt72o+t0IizJNALjqirj6kWxpb8I6i
K9KHAIavWyNzVKLg0kcKGrrPCRcoz2IY7xjoAECKrw63xUUNjYGqXCAVEJPuIzb7
3lP1LSxOdRatntHPYb+qEyPdzDHGgHtp6Lz8zz9Lp1mGaD/o9f8GD2KFjjUdh5bJ
hSWIL7iD2bso/ogzieY0xv0ioQLxa6GFV0Uk1nmfmrxZ7x9N7JyqMcqUnpgdarN8
KH7O0mRRRIP/CLc4i6yAgENSQKfXXnKCKFTP/TWkdFtbkSKCf6SRfXZsu4cBxOcG
FpGLVe9FB2U45GftoNUlkuLww5Ab1uz5zeJnWElhbBKj0jqFkYfG23w9joz867xH
AK1M+vh6XYCpUFrXma5r7EWBPtOQy8vJNqf4Q50kPTVpZk5fgN59jw8i5oB+Uwbx
kUXvgy5zRxQkpi7kXO4kDSpmw86q0+R/npJWPFY3NXb9bdUlcDvuQFIwOEaoIxhS
ZXp6/XArDsXwQhPzZV1Wi8cuVqwrsPp5qLpg4FiwjewbsbfWtUM3Cd3XenDCagEL
VPsMkQAIb0Dae458nPpiMXa0uWF2Li2Jp+0mGVoOefBvGX3ZDLaHVIGQTkTLI0+E
84hTvD50lWQY8py2/2AjYgFo9a/v96Lg0831RW2LUFj+T855z4e/TwB8vWvXKLTP
+zXBWqbQjfxAh/r/lBghgyUhgrpYZAPrikw3aqWH67v0QsjHuf9vpGjICijjGOZE
rrbYvl64y75M4i+aqVXB3ieD6zrZbMOQ2F/uMkaqPp46tsuMx4he21TmlLe2MTEQ
NvYCM2QzuYUfeLUVx5amcfJqkVNODK5/9TBpNRU16wdOjPPsxB5WRCnZ+MPMgzQQ
//3q1e1rzlewEC9Deymbavckg/mHrgTN3wVD1pL8Pq79F/zV0S6Ec9h3vsFOKgiN
99I1AnQ5ggHWN+4BjhudVqhvpZnK0SOU/iwyy/C5DxXf/N4e0x163nXnVy17BZ7N
MCuqXD5z7HoM2bSRI+H2CkilHgoJH5t7wW+M4CoCvUftATiO807vNRXtMV2CaDsj
BS3FSatMdTaeV7uVU/K5S9boNegIv9dB4MA89fG/uIJpLGetHIzv4TNp5kWR7+Cn
vPL651rNbc2B0D+y/uRaMX5NIwu68ycA7i10biBao/c6cF776HhhEFhezGMRmcX3
riIed4PN8j0v4aRrTUQOPHVfBIGldn49OAGKFbh3dPl2YW7KnKF1lxzOa6CPUCjh
W6P/ex2vwwDvvgkwi7AiwzWUaDt3lQF9odT23qc9EvS57OtDn3CXR9OSdJLK1R5H
A5qk6e+p4qExwtXIsapoGek2uPu57oCSixST2F8EkI4kSgqxosNmt4CsotiMGz8W
kpiYAyBifDCxHmjqdvExcx8WVzmIzIDDG+w5R1B1tARJqQyOznfFDaK/2ay8/dTe
1g8cj3wPKhguB+Rn1ZUCgWqromlWukAFgvud0h/inN6lCoHV8x98I5BHgjD9qLoJ
/grkkQ7fzB9LKAF3I94eoAI8IJnosIYJW+NQdJSGXFFct60uASkINS+jqq4cUdPe
VNMgpPhn0CoQpNzjd9+BGA9jdL/DqSox3Pz8GKo0NVYTMqNTG5jJBvYKqFrnUpVw
6hBNwwIC6YlxpVuKIo/8X9cpQnUVgo7makc1JtoPBm8P9PPrT6blvETBqoUrgJb8
a4wUorEMbFYY8p81wm42wEc+Vk0inyOJEEYwGV6K00sQYy4mbE0d9basGDup5DP9
lmaiV+N84isp+YQGjZDlwjvRLEPyZldlWfYYcbhE27zIlnCTA0Gebn2JLVBvSEXz
t4Kf5S7wwEpHOiL28/q9pLn+V1WeR4f5wmURDwnceEATF8DMH4tl8zRqbVi5y7nk
kfVZH3TA1VEhXCsUi5y17xWdZpa6LZ/+XsNNrUFMybc/uULVt8gv67HXXCu+gGF9
a4PDwLxZZh/UeejHPEc+vMqPf8sCKRJzlA/hoyy1SDpiydU3I+tZRRH/uylxtMiH
3eZRqBBkTJsrD0STw47YqDjBBLQ6Haxoh5aTKTpSiH/Ofv18TyU+XA3vT3ssI+DD
IrMNolrwhyyAOPvV76W+AGNKxKq9INH9lhRDlOshG6tUVYO+55nXmwPA8inFVI5f
T27idmU/1Tcesr6emJCRfAZUJ9rGkDeMH8Bl3CoFWclL54K/vnuGRi4Kx88VUAkK
dhVUQBiT3GOiMVJ5t2tkLyn85t83wOVYCooDa4tVlOCgznBZZXSNBQcapoZ77FRu
3OYvEnMimrn9JIxseMnJI5aQZMXXGIROKg1VZGhDyaMp9TxaG+HIgr0d2mSaxSBt
gsOnBeIB5CjGI9fj25HIFsMvBlYQ5UsrPa7RdlT8QEeOnDitk7HFzpvCS5XFZGGl
YHGUgplc3C8W8Gk1l24ubt3CYF+yFbkU6kQSTfC4U1vnJN4rinIQcigp1kX+QATp
j9oA9icjIs/7ixkJVSwy4Gg928nMZpiH5fBIFD4rXsF0SICg7LKGNTS0r+kroW+q
bqt7almLf8iFPV6/OOnpgZ3LrJY1wXHf0KoauD7m5VbfJk/s4Yp2zmdeOG+kN7ee
2+LcJE612SXVnEMURO7gvISC40MhmVFspBvty9nGUsXT472sj0O+NKsPZhMeqlSg
4ltCy/pr65QPdrtBcPcvAGY4PKphTVLlICWg5C+AKlgwWVYdxwWCaRtxmr4IhuJb
sjx7+CfxbYJhTgkbIbjKEt0vqvqmKBKOJ4trCu06AuTJsoaqGHwQAWjUJ6vVl5Dv
U1mIjBWIc/uiBSTmkm88OQinfg1Rsf9gu2ahS21Me4wOD1Gvx7UCJZJney0NF3/h
yF88DNw3EPH6tKQwJr9Veu74TyKeb8fkzXGzme7CJX0uSnNqO9sk0pQ/JaIobWvr
tekKYfNs4j9UtT8QBy53BPmX1Bto/cZD3gsuO4wUuTtBj0RAeeLwDTGX4ZpkJKBq
rc4Llv2nbfN902eDWOA4+BMND4Vv8Ato093wY4IhGRYebAABgdmk8yInAYmvdQhO
RKtthaqmbPIE+udfgRWyA2yONZqvd8dXzVKek9j7O6OHVAMFG++YXYill7SHh7CW
wbpa2kDwXs1IAGrvQYoKwCdi97F+3W7sf5MlnRJe4WtliROkeVPIK8d3MgOg5TjP
b5jQEJ8+oP/MtOLNt0DtPgbTVBfhUwFAavXx32dMErp8HHVLXxGpXtBmC5GRiaTI
9kVnis8kLxscgb7KAIhkasF5goKkQMiCLQ7qOj1zDSMeyCiBaQWjjwmCR7Ryj/RX
81UQL9BPY73QXrJYojmjybq3HsYvT4tKsrTugvwydX5L0PX7yIuebpotBm3U56IM
vJtCDYoQzMWY+3o1X9I4bwIeAbjVol8nySfzOZBWMUAKD+KO/0hS9JBN5CmBo+Ks
wBykTPhAdtLtUaLPvaq/7OKuQFMsb4a2jGHxCY6TjYLz+TmtJRYwt3t3OvQ2lmYn
KUYK7p8eAFX3yWOKhFsMU9elWY0YTetQfKkHuNB1fP2jqV9QxyJkwwDVAHuOKBue
Ta8Iju5Mwpt6c7L/Y0uIqQP4ziwsTvi1m37K+ILS2dJGqRU8Erb1pE9pommIeJEx
ZUUOa5vIqaMZlq8DHAL/1dgOpaMoDtIu+/oUAklIpRB2eeOVS3fty3LlFK05iXvi
s/orWp2036h3cY/c1w7IvwwBGNm7KMtsnANDHwwxbsY1PBgTrWFk4fjH4nrPNW7Q
TDwxDMajCC0YNya0llRxek6D+BAXeXW8S5KQwq+wtetfDtlASjUvc7Nb43M5h+K0
3K7DdXZxlPKJK+l+CTNuLBBpbaZ44FXPcHeQqc0rYU94QKNZip6YOB43vY4a4ZrK
STJzq1GhCfz/Qwx+/4/pYNZPFr8WyP96lt0X3aRLZ+fGK8IjC0T4wkabF0yDq1C2
V7tP3oV/cCjpca0w4NCA3yk4F2HSB9P2BXR2f2ketDVHJpwre8+CinRgVfGeZVyQ
pFVZvlcJUrPwOT9A+9jOdjxXnzzpzse32O1amMs99gOXHWKm+ywaXOb2sdBbbOUD
jZMc1RjfVWePIavvM46sx8XBp26fUp3nRz1NLnDfsXxbEleoi2dtb0hNGlKHlYxC
BgZ6u+h4OzTq5FIwRIGEWjspjH6hSK+MY58kso+VxFlA0CGyTpEw8ldP2uA68wGF
idySgOZsS9+UxIG/0XncA06LiJpaU+5Kkew9GnS7cHZxyLV1vRQApCSsb/qOTp12
yvB8kYxewV7tOQSuCSp8Q3AgYIGeEf0jqxmwNjb29ZxRSlfpPblzewY/dTeBkXJ8
935IHbQ9yXLW87RBkxHq1TjKyWcy0rYySyDAR73AkX579+9i285rrCaHYX3ynS+d
FFIdwkhBhIqV4pm7vV0cPrASkwt+GnX3KftBLQ7Ei3KSR6vmLWEehyAEmFPBxU8B
AiABaauraGKdOTMte2yx6JJf58p+v15nqB4iUZkkXlqACvFv8yL8kTYqUI90UYl9
L6lp9puyZwk8Xv7PNuVT5YYrjmco+DPF1dZOqJJ2awtLpk3tWi7RyzVsiP52vzRD
P9E4DjbEybRJNFK/8Gh+QWc2+Pn9MH+4iEK7YuUyy8f3B4ljG/YnMfUB6Wu6Q1vR
85UE6U6zhEtVenSE9lUH113z6Q+V0lK99eFj9GsoJlsn67AQiu+YD38x6BoDiDTh
SmnezO4+XHdcOeo90ILqwF9vzzxf8ReAuCCfq4KjXtkKRrJeXOBj+6VQFQXZ14Kf
LLQuLeb+sZSylp4+OaBDB0XhDPRiKvp7AltBlzebnDfOYfIzvKyGsFjZMKJZeIyG
rqbLk6+tgf6yN94e3B3bHpWe98B011X/QIsdCn0b3koz1GJqDeenosd0rZMmdOAD
IIcMePjIDvG+1WviF0/BXRnnKzcdcoXFAmBKThAdKxdLtbI7s1uytMAS8jt2WmWR
68Uf259jmgCGPrSDnjsGSv8zTIQ0jGQDjzQ0c7Bshzn9cneWc4fFMM/mrrurclql
JW0ELt8e+W/UQ+vx2NNt8JTqbfuCgbe41Txryk0U8UXnKxpGteABpfpaHd3h6H/O
5derOEelDdOKfay/52ydhSp0Bf8EMoGJFIMn/3eq1k6+YTkelc8vOaPjBQ+PkEvX
dXydCNQ1JHcd3rSYa4R47nqnJnWiit3SP8BRqo9kafbtiM7mraXDdx2/n8ZUTsax
JakI0WFtgnOCqqPj9+Qqh851DAa4D08um3w0Ouk5l9/ICj1SIrzv8KbhaQvTfLqi
XdS7bTbi1KK9e+ZKxsiKcKT4gkGbK8tYia2IMlUVsPXVWQsXhI/P+0lP1jhPo91V
KJJFv2P+D4OreZ0Y9Vdz7cHwtC8q5gLUGvAmJ/GT+OC86if0+OxkgCFBue5xjMdh
HdDn1wr79vKH3i9GcbiW7DR8lMxuYf+ujFQNqEsFadVvKfw71SLWs22CzL+tmWdL
PcSgHkOhwku5Q+VLkoslsumNVfPYZ2Ebo3NWky3WRWnVNgCeQqjBh6LQcKGWxR02
fwDyosufRgXQRUrvz53aeFiP0IqftYmX2pE2pYCOsxPzIh4w+rYy6UYZCgIr+ijA
gCVY0KjSMmoIXtjg0HD/pLMsSamIlHf60O9zsiqgOdCsXqp3AAdMTffsKfymV1fK
pSRC6gHgUAWZI0HGdPJPp/WZDdJW4Y/h7adAo0FQ6KAgF7PfD9PEoGtjwVcEn2qI
7+rlJ7TMXP73QaFBxNhMDJiMAlxEuhj9XyiuYL+J3OnMSeWSP868kq+dnhw4THqs
rEPn84jcCz5fLy8mQGg7YtIyV7uI88UDQRY3rW7XXQASFlp9PDPQlcPjDDrMtUW5
+qC4mjnm3Nl70FfW8OX0EpIhDRdN+TC2H9svpwgDgm0zCZCZscVMwP9eh/PxYvIM
OEnsYGlFL5IsI7rZ+zQLu8NjYMnn3iOozYxMFhVsS0IOhHBRGyofXWko9pLzZuUd
muIg1JS0jEGK7H5yrcMMfsR3KFtyLwqldHJ2i/KWMKBDhYmYUc+xCUNWPyDRQyu5
PDfLqkmYNivXrmmyUUdx/sXQyhR5Sxu8F0ODk+g0GTaj8zbtkWvnHWLDLhQUSY0d
hYYnumiXedLiehX/rPg3112pXINra13oUzIZz4VIDhIDmvk1LiAbtQ3B11avGgoH
w9XyVVglolsjB9pKXHn4LUgCuX5cb0Tquvj9zuwe+uSRiAmk2jUEgz9JsTp+Gp3C
9yMjb7A/oEPEjUPnVWgwLOkdb7b0QWZASXJNlaM3RyVTo4qukK4PkuvTKw9j32Zw
awHNOxrF2Vlqi+SSByWrJso2UMQRloSeaL49+uy4hBH1qyQ4U54X+qf5xMsQhmzG
XktMDvI/qOIIybXgLn/1Eu1pAjzQHWFaIK9PtrG6O+epmQYD3Bvt4U5vLMLMbeki
6b8VsbDQCm589FEdbv4le2F8SsZOMNsTMhQloiHPz/pC/yATpnw+Ybj4tCclSLw9
hRZmeASXhlb+bBbVnjDbUh2e9EiqPwYv4xYzJlZsS4T3D4N3FFATlQeqWCvxNl1f
fpUBsGPjI41tTJZ6eREeOZhztM6+922UccQV4srUdu617YYFBg3MZ3Mfbc0Dr1Oi
rtce347cHWCEVKEyT0DuruvbIZ12RcYmYOf98BbWC7w5ok8+3yMPt+vGpHTFF7j5
UfUyrElp6uxzRdNw/MLHfw2bvFn07rrOita6b1TavxS4EnNfumhgfwGdPUxAVUHJ
uPcf98xK++IOP+Bd0TAXbC4us9h4jj4UlSDdUBWXYQ6Fzigw8YrV95VrOdjY50vF
V8rJZkAYobwYbHvyhj5IlOVcwo70cLOhkY/Jw8p0cH2j/5F1VCpPKpjlgj+/rIo4
O+nzCZnwLTJD9uwgJRrA7JY/IlAqxrSs0ocgiI4zbOBB/shod+VCY87KxA1DOePk
Bn5H9A0owlc6JWmdPI46JPaQHD3ui0GBYRKbVIv4JvS8+ljLqP/JQDk2J/vfu/cb
z+h4isc/ghFdxumc0dPNvgv9uuF2cTkpbd6XIFmV7Pt1UDwiZRojvw2d8EzplC73
dec9MsOE8VUJgSBgRd+AuzL/1qly+XT8LBU6WDe0aZlRfs2hFem7O92yVszuB1Xi
7XRuZSSN5arbr5YGwj7Uy7EgYc4VVXGrwesE0TMe84N6OvZtRdq75t59owxhLFWa
MdL0y7C/acZfBOVO1zM6onlPDOEnXxO1C48nXH1vBYdBQkiLcr3ddwhb86NVOP7U
zCTayltOGtRxjxser1AT/b1Z4hkU60OqrfyoZvvuGev0D1hvqaM7OIT/kMwTem+Q
13D9rSiP1rMmuNWFkQ1Vw3KfORNU3e+G9StvJ4FRY+XjkVi2Gr3pB4Ext4VpERnU
gmRH+UYhK/AoFsBQFpq1pp77KiXjRl7b4fM1DGSm+Y7989UJMs4zSX4O5aQnv7k9
OuPIlrWftbF4eocWwW7cZSfd/Xeq+OTJ4vkHZyEXJefm543TIzDGkemad+GRf+xO
CemWci7KAeot8EemhZ3XAivi2nJ/Ye21N+pb5XOtjCTr5BpOLyTAzGRy42HXFcQ+
4u0+CHR8HuF41fp/BgE8MAPFtTxGV7MqjHHuuSkwBiR2Gl6Oth6GcB8U3o83qhvA
+3jMvTlvQLqTevgzvkBwMDU5ZlqwY5vdeKrjF/uF34m9p2+zksZ6FTY+0VTbKhPd
aDjm1zqwsMWT0OIQXgWF5rHhzZbz/3ZNY1WaHEOBChtLOcVuChFPbjMmJ9gOHR7l
HOUWpruA6MLNcdyiNiwzsPXI4y590mIQ8gJvEJHiFviXKpPH16h7bIpB1iX0x/VP
3rgT1BFTYptH7936JKA6N04ZBNOzLtKTvdtuc57EK/P64YRcLURh9cLBw8c1MOqU
aDeoSSU5MnYsv+CwS6zPN+NYw4s0Ysb39I5c+v+nYjla/y4yWjF+nC+lodbLlAAB
xH26/tg81+TRXlrhJQ2yZwLKD8E8eDGkJRteyEQrZ6qLXEYDedc2kb0vCTIziSW1
zZIhnMk87IYt0BgOz+tvhiES0/5zd3TSJfGoXgFsjvSqRvpSDL6vSkf+CG3UsU/G
YkpCn+lpWBV7gyd1qvdk3mkRLAQ/ZrFk+Y+PcqwdFwvne2Dhzg0JFnZ1bhIru/Nv
FOn441nEv69IXkT2TLtR2YNj8vhyb2HWkxIrrAChXgpo/w59NpkFElzZcDv/DZkv
AZJrQ7rTtl6eYDZrSdPaF6xW7oAfLbWlKpX8jZhDmBJ8Koezg/wyvFmGxrJu5obH
AreAeBRB0wqQ7r7wWB/iplx5LAStVIvcZFSLXKMVxl8ZT9D2kIQF6AfnFbg8QY1F
0fv9L3DRskGolOMMEn6j8S4s0t410+cdgO2/Ry3ZGUN01P67zHwhJMnJn4Nq+1sQ
e45OUB3Qhn8x/VFbrQC2C1nDdZGyzHKT0BlnUOafDv1eIgzqxoOCgzCyxuaHZdYA
2Md7TbaDyLTiFhHZoRWa7651Lv1wyH/8NtlsO7CJnpxBILayi9lqegba+0C3JtGL
DQsqEHZz8tZj/hG6NQaMWisA4J+BRSl4PorVWmt1PkkGqsEmnawizj+6/RbA4ey4
kfJXqrQ4SSAEGjlZ81EeIW9z7FoougHcGX8XwvX9jcZViUnaMzj3TtyZaWxUa3XN
i8xrXUa3iZrG+twUE0D/V1ypr+x8/NcCLGxRwtXjb7+dAoBUPqaBIdfftF1Ah6ak
07V9k8sZ+L8USSgSrZA/tPGfSoBytNeeV7t12QFQmXI3MnJtAQUtgcdOtEb46l79
Bw3SmJFvgQJLVcgDqWhPlf3ofPqw9pynku9bQxQIv+kjruC1NfdoVxyVSh5VZQH4
ITnKojX3/fri9GEkMcI6KKkvynigLOqtw+8XyrS/0WmnxsKOYX1ZqWR7SwDA+T4j
2rhmUFhf6ECeiugfXuldoUg3sgJQSrrMasa+IxIUYQoZbTe5AsgQajcZEq1YInR7
rD4dA1xVoyMG3Ojaja62VyDMy066RlP43QnY55gJzZ9TQmAwmyAoAPXu9ih4cf/M
i9LKSSmg+BA8WElv0RNYguqg8WHDCke3urfnkRqMoAVojSdgQYye6r39t8utzuOw
IVlTb2KMeh5FCTf6CiyhyJLkDpIkX5mJqNYjdC4R9vHajIZ/4NIKpSfIuwCCcwfZ
RrPXgTGZ6OgE00lyZPAlVDDNqzjcAra48FXKNacbMp+JjkO4d/BRvZnXuCd/8oQt
YiM/kmCswazLU1AELrvLyFqAR6YATzhlxwe/56QRX5LA9Bd+spb/cpD40+ojLqJk
IVm9Eh8YanAHy4ixUGU5O7K9IukNOz/kHmMTa90YT5JQsp/IOgCpK3nKBWvg00M0
+fd6Hme5SHVLu0wUsXuDkzIjdJW+IAfcGoFn5yXy9SUHo3ghApfrVsqZ3v75mz5l
pNdB+w+h5PKAXno/RnzHkHQJcUdm48M0B1TPx0AuocYTkEytEduwmyWrsMjInANz
kWhLxiIyi1gG3b7CzxV24C6WMQ6UB3S8CtI6UL4AuV1yIibis/MWtuqG4F9WTd/U
uopPH09buOY2lYAjRKCdatO/gYNx2J54MBxPG3G6/11kkbAAQW2ju9jCIdYz2TU9
N3pB+WXp+knIke9pxuR7n8dfmJgHbSHjb3w6Z3bvVzs0qwGgrYNyXSuDofxs1qW2
FkaFg7NAlvApRFiM/+UQP1kqZ2YOBe1twXJs2G0mkmi8ActLTTQ92nNX9bLG+Tkv
C0dgB60qB/shGb4xtZqZIVHPlalgn/4vkWbTZLxwmwnPFGhxEfIcGQQVVHoGMUgG
4g+MXIWddU0Dm/5/eXz6OFRu2+HCOm39lT7vEKjhZ2iCs8AnKpnrn2whKUxkLPSp
K7ZuktwXnuQYkh1+VAa2XQbr50pKUMOGF3On9JxUUr/P0i14ntbvzF1+xcFxserL
qzSRfmD6BUZ/yPoyJb9fRj8/cKUFXjFYm2O1Ta21HYa+/WYY0pwhl68gIqQbjYRv
0/zdnlrXc8LEIEJ4dy16UHXa4epbDAHZQTMGvReT4R+Rj2Z6WUf/YUmnKErDDEYr
ambO6NQ0hOhDrUAAKQhsxpqJLKYk8nmfbyuEvrFiMbzRSLAXJSngPUEmP/JFjA5h
YKSHVTtjK8MEiiB2zScqRLFw6hZsqsap0O/GiVvZwwjL9j7frgdda4PfV34ieotW
q4T86ZLZVOcoVQMzpEQIUx1n/4HLl0QhOv5FrYUjfaytbA1Rj5HarQZZte9dq8kG
e0tH7aajOyWxdj78fydfsNP4IFTZxgG/rc2sTLnR534P7lfpkMxhhyUiZOOLMVJz
l2GYkBu1RrXBzEtdGcvXV7mQT1UDgSZUTlbDNXmI8RjqNBLKUysBEabqN2z7nugW
95xCJF1RZNLVtEsHpevZhKeGez533sSEFzSbSkczjqQ2LdLZQRgx72nKPCPdMEq/
rpm8crScFPHRKYHotwOZ7bgBKQUppTXE07Z9PjIJOseZ6kK13rk2MoTiJfNDXrEX
nyUsZmnhejX40SezXXgmw0dn+e0PYUJRvBqUyoE/14sfrktaFwBGdQS/YU9a3HB+
I1GYkBwAc0luqxIUFovwLvyCQKtOLoV5UlqcEkzuqyEjgkwvlvDVFvfe4o6iDIag
IBgViycMpSvRJW8K5sObIc0Oqduot0ebbS66lUIGkuGAiwgc22ghvSs3UY7btU2k
EtjRjt3uGEQxc4qKOtX3jgzdKZSKZodYL8CbcOHEGdt2fU5YzEpbMe+uoPapwczf
2/TW9TW+9XjoTdG1OtdUksqd50ma6xggapGqLMQv1jYZL4cFPypvmGcyXupaK0H9
edGTwo6Nx3Axn3kAq3ZxUhlYJ/Gek4xeMw023LiHRoPEWPHjQ4/lVbZ9R1OExbUn
JyaFxUVKLii69Y4+b1nUJDr66rk4cSAEtPUdt4yg0TiYDPCZuiS4pFF2KZK7z1A0
jVLQFOY97Hm1Q3ODWCENefm/I338TJOm30zhK/qkwj45APiEXzZh8Y8Srav8ujqS
3nm8bmTzxbBND4Fv9f4cx2q3prY8yx9sLzMpyqzdN5PjP9I9fDu1PTOW7eELYOCw
WrSbA2dIj4F2daP2npSMCyF5pd4y4l1TkFKLs+ivTLBZDkkQxYsTI+eSiWSCLBT8
pgkm0vMwlPTtwWlvy1SHBUmMegT9B2E+FZw1a4zZboT2Jj3eDVc+kb0GEdQQdm//
gliPHPcZzSvLC3NylGoRoFkoaOHHNtINkAS8tNYGmnNIc7I29bBqLNUlM7Kg6XFM
952i7HrEiR9drt9DiHVycVT0cbjV8aNhMHOip9Loyl8DwMLCNO5gipnRugDzR6gV
RR7T0/IZE6H5CuvwiUkIIXP6nV7AUYQioSgdVWclBVJxsBXLFsD8ADpxLexhjY0y
VPWQNW47QMR3nBupE86tfxXjckuruEE2zS48sq9xqUqX5egTryrguZ8An7Kzg/Ua
MLst5+1EOWsHENDQRl5aB1qAY765hGyJZQ/gW9IYSp7sMTn+UAsj+8n/bD5mQZnB
JylkmJXVRwH3fzOMdGtLPg+h+bZN5BOcU3n/Lqiev5TF1KNO4gxMptk+mTMOL+SZ
IuhuTQAEkL+SFeidRxOmwOeg7Ew2N+uH8sHEKYB5p6/bQuFlU1nhF94wkeImRhDt
qnvS5lhuV2e7xerjI0sWU3D2p3xvYxVk4zYyTcXMyclowCCPJXPOLWCMV8N+G0l3
7w770O8PWJFAk4c5D1iJmC6c3WgWiSAFBKvoY7F1ILUoqlz+Z9zvXkTM6acEFcHe
ULsL4vT+D+N4grzz/3LGH+lWcXbk1RVbkBM663yD5hEgAi2y3Q4i+8xe3uYov3f7
+Ia6/3dZj1Ll7/TIVl9b6IoMEQpi0IBYKRY/kJKZimti6FYWjhIffdwdE3j5eM0d
sMzJxnXFf/0Kna4TdI0tywDrrCCPVke83TEA5AE0MLTT1Jvq4em4jno1oXOeq3sB
1mgNYZOZaNWJ4bQ5yjgmRnCtTlww3KXNjVKakwCt7Ia4xa8po29deTPwNgpsTFte
Dn8GEDIY2T7GFGRm6ldBGySoeko/cm3fbUpJ/xUplmW8oUy4TV/jCuse0AYkeUSz
gyx97zUOFO7kzFswL451iJkWlmmlaND8pAiNXafAtb2n2YS5YpVmVYsW0c5CXN3m
WLQ6r10SkecbYIY+R+4zt9vYb6aYkBpnkCME6EQAA6G/QEGjKFO0HuRq1J/IhHyX
vSk76eFnmvl+UFk/vQMZPs0cyjwHyH7q6bzDEZMmDVqqYjx1X5+sNC1omjXJixVe
oupi7m7NC8q2yt9N3l5J2Py2T5oiTnX0HZdcDl9M8BKM3Fzl8P7EPf0KDOt7Eu+v
2Kg7QzBXfcDQgJyETvfqzUTD9sOLJ+IJNZ6uVWFJyT+jceS/oTyPiej/fkv3ISEr
QgYKNeBU1w70tscW2wDtq+PCv25SgJets9oapveCiRu3nxUbHWYo8BvdjBAeSfsP
B8URrArLukdvvKm070lESUrTm1joJi9KnbWHpBYuwTdjcYhWFUnWfzc7vY7zP6lf
lyKaEqaC/UeOsmRm62S5lgV6l4cE6aIHj6XOlj4UWuOnVHxakpRddZ21vl1rpe/a
xEyEwfkNQ6jCCBK8SV4WkvlqcTw7Bj0ER3PYE3/fyoI8ylt0++U9I5gGxLMzjsyh
oDteAhtGRYyA6PFaVkQrriXIyUeZuuJ49W79r0tIJTC/yl9fl9Z+jodJVFtsTyma
ArZ9apF7m2GfcY1FyRL8ZkfxOh1Kv6//ZSAhX46sdbzB1g01S81RNHvRmKKUK6AK
xBvoNRmzy/popsKOA/zZ4qaiZof3XJK5m6jTcX9uTdCEfPRat+tbMooDM1JqEsox
ZaR8dd0A5nIahat9vDog+mTDMeBpOKu2tNPV29sVRS9OnGFvXTW4aMOmx/qFne/J
8g3c8cjRdO3m9aDOYD9HfNa5LBE2rIjmTROdi5MBXG75RQsSD0MmU3bT93HYx6V+
mKWESlepL45+lkqIm3owm4LspXNy3mlyXDIT0Erm50IhMy/2IMcsqBSmlM/IcllG
ywK8Tfqq041zoa/484BCVtVsSKUkPI2GWztnANJny877G4pVsrxBTW+gwNuYmrs/
m2m6NtiUBhNQgsxTmHT5GqJJqZt6wjuEw1nhLV8ILmJG+uto/2li02yNotnEYXF7
Zb7kSZ9YufDev/brh/KLBteFRE1Kg6guyTJSFGzzg4aoTo/Ewr9rSkNXMcKEfBCw
tG5G54gIOIL+EZUabL0HQMLgIt+t5ho/91BRTt+J+r+PVb31XZU/SoX2efkExcKW
c/ObiCsySn1VBdAwLj4F/eCUDBq1EO4BAEA+vqeI/Navr4kVQ2zXpZaOR+2AogQZ
rSKxCG/W0lKxBNW2zqC+Kf00+YtDCSGZZ900es0vp3etNSLkEB5LfEWUYgRdw5EI
KyIwcCiN3Klf3TQM6PGoPTbn8bIhMbrI7J40dFfOmPh4VTXd4BFeN6nnk0DQxEjX
Co1woThhh9QUmdqHCIZ99L46YIVHz5xlS0QC7QMcPqOKTdheiSh6CXldc75qBNEU
58vvp9goxWIIcCWTOX33ePivymUBnD2MwWLr9A3pEJNyGbmc2EDC2n5/o1yuN3gV
dK2RUXyOZ1Hxy3kGEDW1UlLQfpMhQFEs31Q212APkDC963Rj9JOPCc1aWiQNo9jn
IoN1WOR0q0wjjFzog7gD+OaYN5lID7UrZzm5jAumyB+oSemYba01BTz/iDQZ2o6U
k9/haiD3VvLofLWUtHFEqC03y3dAKGLOcPkTpofBhFhuzfj/WVZoklXht/AvC1St
bH86/42t47DM9jgwY0kt6VyiWwXCjjlue8+7Ygptl88uC6DvrNmwQ6D4jYNYNgzj
Wwv0fyMU0Cvnh8mSLmiaSAS9DAl0A2AyI+HYxJLde6lu9LzAwJNr+B9BRPOKdhkq
AvS9xlFL3hbSaevY+jN9gO/Yk0sw1fbAs9vTApBOuLd1Vpv4Gk0hW52aoTGYFizK
38J5Z3gNiMCjXPB3isXmHZLuuu8aF9FhL2DA9C7d/jVVyp241smsfTXAbAhV++e1
bMgSqG/vaPeCThMKJYcp9ClGhahTiW/ogMc06fXQUSriGTIcOmyc+h+TDPSGkhBN
jGI2wSkeuyI62wW9re+U5unJkv9/SpYSHKRgyxZeLK6Nfi62hV7bZQS+nh/KiQPp
67r+3fkRWJX6aRJHM3/VtuPd9FG/OC4D19sYJFQI/muqDvcyoEVpajvBDzW5AYlI
3L3/roJZql8MxkJVWeZaj/4RyFfBfVBPuXLX0NTiGyheDK0o71l6FosoGUGKDO1Z
of2qaVN7uUs89WcNP6PNU9P5e90yhGgx84PDC8j2GVwTatakzLsXOX5vUwFyDBAD
3N/ht4B2Gg6AslT9UofavtZOCDun6HTUEu4Xf9kk+Zf15QiXenpvJxYv8YqL8v3Q
DxWpJrp3ISCbxZ+RjxsajSuK3NaXy8bmAewhkReNB3Er2zzeacSZ3FDJfIofuAUJ
CsiJX0QlNhC5OSSAIZZo40OnGvB+elerfm8mcNIEjS4PlZrtnanlv+NsikxRg1xp
ImVWBlP3JDYk3KrCArqD0rsIgKwrv3rPuIN6LP4MbkMF4cdoSNgfH1GDpo9tfXlY
KvcvmnLiMn4Qi/J0vfKgg/tONOkriNgRHIM874kGEQvsILbUCDxw9rDOwRDzTcRf
CskMFlj/8rUT1GvmjKd7FuffJdpUdQJlU3e9wtilZ8N9VGDfRavZI4wimiAPruMV
V3xUnmlzPAEM0H3K8E7tfd0f4pCyFfjvVyqc3eFXPWJXWxblthqAhDUIu+SDKpSn
SOIJo7wpUlrMLkCd89Y9RTeDA+tdDKX9XOWSuS2h8m5NbuY6nbE8Qv+se8GT3FX8
ZpMTiWnpLUPaMMIgX7JL7EMzp2+FeoYnWEn99m9WAiTzEy0hpvR04pDFdsXNuCwm
63/aZpp7Cpk7DQWPNKZbSRB2Cu78RFdkebZm5EtdkpC4gyiqNH0+kle2dt/Unod3
MmTtdBqdz5nEiRoo1KmtpvqMwFetlaUg2+VTu1/zBUqITAPmkFKRuyZjdoRi25D8
GQczIoouYPH1O9lDVhdXbYuFk6kWLWl9mDtfZninAD55umAJznGOhgBGOslWy3aQ
h5PpnhL0Xg7WhiKg0/LtdztlgisW9fX7c1CueEp2iImKxWhbAwd3/TPFDADRAr7N
UiuTsy0vlOvDlooiYtkhsuLkb00I+BBq1mdCEdRlz7ONQyD/geC9xVL12cPapNtl
+mi2bY/03Khdmxd0eL4yRihSKb49FcVUDg3uYDAuV5eN7fxfSVVGoqsTKcafqond
RifduXXrdDhw4q5M8CTxYN2lTcaA78d9UFFy2aX71japNY1TfD0bCVsKnKFzchVh
nyhYGOzjd65GRbDmp1Wty2MPFSJ2WuTWmqjH/jwBLqxJfC0otEx37RvAH5RibBdv
fwsBV1+ndsGIWB5gn28PNANhNRUZ8LpcTI5KR2fdxOuNPd1xDB614VudYDVydW8S
SZmKLFl53vKIDV33FV4oYbJobdn1VJTAeuZ4TULWQJP6Tg2sq00RraZgO/461LDU
dEBCsr9xAcXVxJXBDfw3GjeXBnFC4maP2BkTtMe1/YoAPJkqB+CwF7nXocfFJgiI
al8RExmeIYuksQlIWKSa+a972V/6M24984eehldcPwOJGRqXXZIj20vazqG/7PEk
hoXhGUiYy/r9IRs81OH13FFPOgd+hf4TzBBUvVoMWC/2ITC82y0lRhoOlRh1mFxF
+lF+9hZNjFDILllTiLOp3UFQ0Z7D3oREGQAOw484GVDqdXXg0aXCg30kTpqVClt7
Fur1+R2r8A1vAaksb/j0yo+FlsLuYmvwxyo+QsUqD57Q2ExUFFDoWtFR4oUKMyYI
zZojkVldjT2+Qtj2UT1l6GzUhwz8MSuuqf5Ud2ZdERrIK0UGV6SBlt1oESkeBBfL
8t1dx7G3ge/mhe3xfC8Ux7FFfADOullXRQ7JXDk8K2ZdkOy34cj4ckJeHDoZHVfC
zdddel1g5gLcpCAS82WSRkW858u7RtKydKtTlWlLLSvY8wrLIvg0fhqbLBf2CBYk
lHUlEssPHMBly3Wig0ZgTJH9IiLwZztui9OA4np3idljcd441Sp/JaKLVb8eDqol
60pKVccR1AgHCV2zB1qX49NZPSgridIf24D5gVu/WlYW6wiWS8u9kZji5VA/nlKY
jMVgPLjOL2KqlSAo6u3C8MUvLltIpCiQiycyQFPNt6TkSRJcF3C7RgDH2HRqerAh
TJhBI++cVvqqrQpyD0V/OAF3vWPLXNlIh6IxpjPEhdPKWeIsNS723m8dv3sSw+c4
BrOJG9V4XJJ+xaps25XUhE/Ns1CvWjttkAdk7xytJNXvT7f+3KJ6/3tNSRUBpiWc
Te3CY3tcw2I3y1qno0l/mpfPl3Lh7BMMIxR4F34JhKgKDjLgNVpvGxuxvz3JwvDW
/lqrncMqAVPuON6Lzor31c3f424cY3AEkhNOa7/XuXnPmw8w9cnaFA8rFHDaJR2k
NIXshCuIJtwOrDaKF3Zo7f4b/tG7ZKJ9fQASdHD6XA3Y76EYhtXIggVsxf0xQs39
0s4GnGwjMoer5t/qKiMm7lvWnpHsSwWaI+mfyPaRzFYmL925PtxPfhwk+22VObCG
RXDsnWY7jL5tqI6vvYwrcNUu/EKZOP4ZxagtegPCFo1KlcOlGIkAcdoKitQLdaka
6PLaiIOVKEPN0sdMEo12NKFl1sVyEJQQ/o4G1jul/JyF6COhJ59d7UlRbBZ6B4b2
c89GMTVKgTzZpLyxpHsigR/aZM3c4TnErLTGNGyYyTRum4copd8AJgrK3T7By+Hk
AytbV5hX8LPl7b9+xPkC0BGoOO3Kj9NxRUmUQGWwbtiEBm+sLzEzFDp+YA1PgHdt
GGuPLA6Iercp6CbN3ywiJtWHCnH627SXwKn1WNxSPTjMdxa3U/yxVDAvchUzVtu8
5HZ+eItmyjvTnEacPuuYkzfvOsW2Ze/vzFNhPkMRDDKEpBKQ8P2R4PHCD9NY7Kgo
FgeeUsZvwaS0xN8HUcaS0XcwQwYFMSTOxP+yYusbpEu88iAAMlq97eD8C4T/0Lfu
Ej4eq4poBdqyDrOrhkZw/Hi8n536vEfaCMQORD/Ym8y3xI75NQZIroiU1NzhrbuJ
W4ppQ00DWf3sVV3Iw5q1qDaJJEXKpcMWrjwx5nD5SxNCwwy0QEioUsGhCw9iyZhH
3mm+jz2eGoI/PnCdHaybxXxvRVbQPv43DDePPb8UgAfGDcbYJ7gHtz5GHINQBH+m
nbin3yK2N/xGVPcUjPUGKk+KHDUf1WKeH7Gr8KTT0JXtOKDeoPzCow8FMkl2I3lw
sDwYzPQ1GcbOWr3nZL0ogsPZVv7WxAQ+H+uZppIyf323kj4GW8hw/V6joLmMtJFT
AHZd4xDvNsbXyw7DPS0JgcAIeYTDo/vjn/sXeONMtE9bzZg/P9xGJx1BT9JYf/8T
Vo32MrNAHLPsv1wXcCKvetEzsRsxNNP7mZ1sp48DPvrn4VLSrHtRJjFW0GKcabbD
gbGEWsWiBGbDZfW/d5NQE8PW27pEjGWwU5EdR80wYCsmTFeQnjQtkAO+0XYIjXq2
dHADxbd+b6oBQQVMqCM9QmmFj0OXP/qRTH/0H9Ci58YVA7uFI0dwuJGdzVKgNXt9
Bnw87RI3rzh2l0RpLuxk1QgPqhGRPI9BRYErAoMnUw2ScktY29eQnNs/fO0wa/dk
mGf8/nv0INRBufEwXPNiNTcngtqikeNFEFy2hDCobIcVfRz0tm6cvruA+OhIG17c
HM5riqjZcWDA9NvIy7S1BAnceE4Sa1MpUGAJL0Kq4bvoriQpelKI3Wzi9ekpV4tK
AAmOLvZmCyLSpbDivq/1ymdfMt4P6iQPqpHe7YXHwSG2ETzVpKEOToNbB9lm3Npk
RjDGjT0tQZanPxiS3XBireTiBA085/Doh+PKzRkaIIzfLFqDLFqyzGxViiI5pDE5
3O84ndQ4NRWOx7TMcrW8wMs8tlPsrdriAXNnZ8VOAR+xhprHsbR+/itKAz5ADfgs
ECgUiO3ZBJLcdr4nN5BKt/TDF3uLV677W+dS2JoTY7TFMKDlK3NKy4QuYuTSzuDP
koYOcbhqaZftJeacsT5CP485HdCWl4Pnr81Al9oThtbQMMtBdRLbEbNAMqO+49V3
GcfRfpdPGJmwmvfOXbN0WmJr7/yXU9Z2jumzkgqf4/DDghTLWAIZ06uLHDoNciw8
NKqsaPqZb6KrXzIwlR9c2wMnEipHYVeQ0ymnSFERqtk1myRD9eOuP7J0HBwFnqwT
RGV4aZKPRPOcyzob4/pukcGX4X/SnkOjtMgLJxZ1sScWfiyW1l/EfBKuzcmtZkxy
AK0Fz0poKXNLUVAWlyMG2c0tR0sfW/XJYbsF6O56SjaYcQ8S0RBIoEarEgi2axgX
/WiAyDADFU4yj1bMEQkh7myZrdL25s6wv6qih138vS5IBCC/Yyn7+EGpxjRvtzgX
8JlXq2xM+8+giV/UkRKauCT9fksfXj/wRJZiFMh17pk2EMEbepAU6ZMQiaI2QKm1
eRuKAUUzTdXIm23OPcF9cQSTsZ9uPmcNlcgwQaZoVaKrbuQt5yNpZLWI5LwHQ+Um
UVG+fLUE9L9PSRSKY3wMZGlSGru3KgDPjudpc1ydXcwB6VB07SIVgjKI67uAPvUS
WN85rlGBRT9MtweyktmhUlIg83cl5Pc1KqSWbj17ZQEClgfG2d3FmiQBDB89Cbb9
QfRhkxaEXXIXWzbIyGMD8KEKC3mgUks1pheYjPts8a/HYaBwuV+/o0oFNP+2p5lr
JGATSPOf0d9XOEqz7gB/fMMBoU7OTYU+NCJV3+D6MkkYK+IGkTyXMbz9uUlK3P2s
0Gr9dtH6ScTuXLRjz6g0W2kHp9ENWr8IvjlSCxYpV9ryLkepuNbCm0riSAL5nMrZ
GCOld62oABoLATrd+AnP2pYuBMXUVFdFd9UekqO7iRZMA5pE2OIouDIh1llDt+06
e1/KatiwIjPrEQv1/DRdYPCM6e8PA3D+WlPtSwqj9nYVTgl3HguBLOhs7nC9v6oB
moODDDuL60v1SEJ+o31t4Qk4TfMEL4oUMWg68NxTya4KWoeZSFXTLNmqSMPxAQci
wQYR9FhLEnV4q0daRHSsNXC8l/H38a1PIKRhTmiREHhmLvNoOcHyXT3tB+vnsI/Y
qhOfpavpzQdIKJuylCbHBAWdjzX6kPxCOQVsBAYIBwu7kjbwQsgFM0omhd/03snJ
DtY9WXhJIsYv+NLwDX1DIN3oxOZMHBKwzCG0/lJQbDf2LPgOUmR77jTmmXjr6k/5
O2+E3vWHMINJiHLWwDHUp+kjM/xlu1AbRIthi6FHN8GU25VvHjd7Psl/BFT/Etyk
HoEqu3YEdBl0gb/e9OdDpr9bOnPpvFfWSs7mIYaXeMAUUG57SEsC06iUy3RqA3nd
ArS+Mn6tH2VyzJptyUEyMhqWWBC0fNFWxthYkF2enl3n1adoauxp0vGktXjSsZa+
/eX2YoAGuwX30Jd/a+ksBcM6+FZ77HhBCN31W62IoVC3Tp7aU8fUXhykM3juUwML
OO0FsBA8iGjqbsesu/Dm3m640K2H87sU0owLXkIgA1YkgPR8b0dNsjfeFfCxg9g0
RP6UOLR4GAejMmYnIv5DDw1f7aj6PDKA7gwyBxQ91VSFRXpdRVPl/E1wb/O9Rad3
7Wz2qjn1i3hMrMqJshYKKayVGBz5OpAF8kOvFQl8AwUSFTTHRC0Zm9eIwJMypY4t
MU83mbhktYt+9qDNOuXcrhPNj3nh3m1rDOpmMbHzni08WKQI9zMv1JDzMIAD0awC
bA2xVY2OKqGHJJkyQfcW07/mdNh6Jam95/rmCM4cbg6NLAmbbhiZeY8OVfxLNSaC
GOAsjC43e6C574g3e48S3mvTQGr8DUIzhLZiQg0IP1PnKUWF5FJlPpoJzxBXhOj/
HKeFyJysQFH38QBx49SAsFgndohvboHOO2QOeSAWa32jcE+eMRSul6YIxQS2/IyP
rJfznUbmsXD0NhL1GHtu3346beM4FhmugSp3K1N9fHxu0c0dVVuJ+vksR0fsFdGT
58rPiKzb1plk7GVlDmYzZpxUypu5R5Uk7mNlg7c2MeElvpLlGh7iygtlzkogA4Cu
s5lKCRELdI69Qf6aAyUpy67XVUu/zpInNIrYZPMkN7pszBANHNduS0C5V4FEC+Fl
Qeh0KgY5yf6mtXHwv34qRwtyUMO0DwzzzGHxNNqduhxlCc4xNv/JIpm59HSMC+GG
JSQW+TMujAxA7zvHvipElSVnjfHxqJno7HwFySmk8GYdesa/GQpCzYu9WxL6QW1b
+PxULaT2VnCLRhBP47H0LRzHzIqBf3lHLK2nJAA8NJm+0TJUlmYPdQlcgQiQjbL8
OTJ5cV0h02I1vliCzO34J+fJ4vHNK5tCKlegOXxwY1WixAcd89dsxLk6+DWp0/Iy
tUrx2IbYoVM2LfJyYMBimeyGdtlIPA6oPTfFsJcP1aJSXSYVUUoJACsegT8Pg5TQ
mKsh4RTgehFt2hrOD6JEvIff5pXOpYyzt8laUTkx7NpJVtcoBqCIZ0/V1/Ejnp/h
0Qtn2a8ttelSl/EHyx3oxnLLC2SwCIJD19l7tSluKaTwnuVTlbXxevm2M6xILEfP
VyJwAI2/Lo3ptwi+yRMX5Aqws30kJn8+3L88awgUrYyP5nbPq7V9D2pnCzIaP1R3
W5zEMCeJYjiyAHEhBFS1HhzY+Sm4KwIsBqbJN6ftViIY3kkUIYRHwMhL5cKGV/2M
5/cHF2ebV5b5Ks0vTZo0iMCayfnWGH5Wy6xXq8iT6kXTwsLvInIrjjdu8iiltoZx
V//C6Ni/2fpoyX7Ylylwrl05B/c0LtoGdzUtFfmJ4lUJl9zAIw6Fm/DliziWAyNR
PkU+QcqJ02qJFUWASYU0OzZRZBib6FaR27vFhOHZBsHPkeryGRn+3VjG2qgH7DLP
OdIodAnnxA3/ZyFlSxCVq4tIGf+A6SujsdG9XBY1BR1jjYUrFu1Wr3H1EMuBZ1fk
GyeDef4dovp44KOxV02hlI2dMTUITh/plXB9b/Khpz9xdPEh6vHkRSPX4AeQRZTl
McCtjUBkskbcMaKIm3K25ek8mMwCVhzJ+yQQW6OWu7pPpmp2Uasc8mKVrbvzSdRE
pGwaZjn5waNPY98Ct5pk+Gn9lWo63TQGn9XBz2TQaR0WcW41eqxYWN8daOBLlUPB
voawqpD3ZHZjJD548jZkcuMpccaan3DUgsDofaZH4LGJhOY5oZ58W6elC6lZmu5d
9Dwh9bwlxWO1oMXv/ipSlF0Ou5LuevTUJuKkVUJoOWUei+jNFgDASxjidWy6hVaK
nubpDYXcUNs85HHxEb/7EJGtwv9Unj/eF44EF6JmDcjACOaFL25gSaXbvjuR1prg
HErszNaHcLX5dBBe+PEbJag5srL9GBFNzAQXM+c117BEj68XmzCRGZATvAmsfk/d
+INhFO1RpjfhejdQ93eqNtC5tsCKOTtfHvhsuPUwNZB8MDyAUXl+43Bjy1FHeyY8
S95x1Ot8gsdg6po1EDgGYtneRIZJOJUFX62rpadajeIaFTDPir1dLkJKyl+Gr0sj
xHSvMiFnrcB6kkhDY3kphwlBZ1xHxbzmoa8mr/aw/WC4XAnJl3JGldmQKafCAWUL
8B41dy1qoYZdxktUanmZb8uoz0nPqXI3F6UIvlizDRALO0TQ0Jyqpqxa7wqznM9n
INEjAnUZvpbJcv1gs+nK0hx0Zr4kd/svWmdrkBTr7ecLIdT2J4ONUmGx11tw1giu
0Em22llaMRXh/uY1J6faOqwJ2f0+hXT5h/FcGNkSXSRhkvC/De7tvQne/NIn8wlP
rlLlgY32WKuxKkkgZ+GWUzbDYxERk/eY3JVU+LGqfszZ5py9P4uJDsK2G49DHOH/
y4R4Oi7yNeyKALtcfshSt6LAq+WXNghbjQ6asJ4J1ldEXUowBQK3hiY+NhOq3K4i
A4wnO5eDgWaIJXPTIispa/OCzc6S+0wVrKb/k7EKjVRGpf/4Qs3J84Ovk8TaZyEm
iOZ21o0aAKD2IpoWWGS6GWeLcUjzwNl2AZV0VKQpz3OxB2FJfZTnVtjR78gEMW61
9RypvwUcI6GPYyItonP0DIbATx/wQ5ocSJhu8Uf207D6eMaPsComM5PqUbAUTND+
hcWVZ7WGcpcG2fQqmb25oWlL5tR9KowF1ti4rE01yD+/NWCwZFbA4+CF6458QsEp
at6+1U+A+QqvfW+XOM7+jwzdd3P2JtDVY3/qAEMoUmKH1n1i72wWK4Y9spQN0bqJ
t6bmT5O5Nf0yfhipC/kP3Iu48Dhgk6PI5exLDSE8inH/eUI/+INvNEg613CvyQej
Oc0/SXLQD4bRNwuRBf3vDMgpHCuBCxB+i/t0CJ/+3iXTywLo/hppNodoiFvu0+eP
LOK/yq2zrTzp16W2QCl8om4s80O4yW6IOhyNEQIY1SC+6z3o0aWgslGadFdn7nae
6xNr4YhVOr+B0QNph+hy1c+kgFbO5AUb2xY3lLFKeFNItEiJHcvRACFqPb94eCnT
ZRoZ8L3BiUNePEzcpbDFAwbThzAadkfjG9bj1dkPLzCYEvecPvQ70rBWYqJ6LWW+
WfbyX61p+OoL17KfwYIPZ4CRisRq27H6ZQCeP9BLR/cMz8602doexWL7CewZhiRO
OyzCWD2N/NDCzXjyAsyEuPcmIHPhrDBZZQt68B9/1lEVELc+RHfpqRyyB35VLtrD
ZCrErC+E0vYOG/yWiwzIljE6EIfZ2O1zMtjW9K3l/FIPHObKPTPqKbJTkRqDU5EK
t0lf7BGXK+Xzg39XBPp2L4jhkib0GcoHtAXT0yl5eNtxiUWyf+LPtToaG0VfPRv7
eTR5ndS1iyt08a1VcPmxadbzWkoZHssl3jsN2zQgvpnwDVE4w4MndKkbGpzjuly7
/6it7n37m7vrKNCs/nCuK4soDXbupY6AiqmZOupjnZPk178wJhAnftamJ6jXSP/3
/d1GFAmNnwC7mReOnlm82kZKihWL3ArwsdmnP1e2/FMX/98fSmgWNM6OULjmZa9Q
BeJfPjtXpTHS50sX54EeYpL8e9h5EWp2LjW8/YMddT0r1JIoAbv+WlQRas5otGhD
071+cWHQoUV9hcIlvhmtaHjGjTJfIgWT9wh0sI79uEE/7D1zf8Xy52awDVqZ/ZvN
aSj1QXYngn8V6WroN32lOcaL9tFm3ShNQgHT4Wy4+En5zv981kdNKFjZoaXmK2yg
PbonV1Uo7CxEnYXCHmkAMvla1ck7Ugm+gIL65Dz6ZLN5vKEfZ1pOnuxWBTNh0phy
fbVTKO/pceK60Q4FjgEWqWzglBGUW1hX26+n/cuaVpuuPwQScCBK/7olBXtgYGrQ
hvM5ACrPs6j1/Tw3V3+9FCnFf939SYAfCX8BWdznvTFNFaorm80ZUHH5tkNK++L2
aM8UuYjlGQDz9zoIM8VQHXDoQUfq10ChpZ1vkAV/5c2dSye+Yvme5gAgGnJF6lqA
ZOqCVr4O8eSeC1YTWFvjrY+a1I3A1rdTWLwDD9SZFDTsM4LnSd4ZtdYI7mjitMru
SMSXIuH5sPEjvYgX9fY3jr8bcQO9zxPF2uPFh9yDDrVR7itlcU9f6pony8SqusYt
FysvSlhLOMW/7VmJdYjKsPPGvlbaYSE+u8WIUNctDcUUXO0/CgqjX2+fh8VbMvo7
d+MoKgEu+YDF6wwca4FCaHOkoXCnUc+5YQC+ITQjEMDNd0q28GLb6beeIZswk3HL
GCaxSBHb9bdELRI/XfgzUzDXnbYwgnzx9eexac2nPa0BxCQG0IXyBD+RU4PuPFFL
W8xUcn+MwxqrF8Uth3fJy1GhQmWfp4C1VwhNaT8u2aqcmAS//0olOyQHPKv2T25j
fX3nkM/D+YyIjJzbA6QhB0lYiyW8U56s5FXL2n1m+DfMjBqpdst0WrCHQK8x5DqB
4qojQz/ZlMxd3h+DS8ATTyHJ3NRbzuIMzLf/IBwAqwkrHlt0d9kx5AxDSCcqphC2
B78qD7/vLVLyJmOd9ETvDNJBtbyy3DXTG1dVWfeV8SCm968UMEtIj6JFoTH5kezj
icG0zH3NCX6/igLOl70jK58CWy9ibIcyXuMwkMmRXBsfvguss+9vzXiWI9QVK+01
8eg3rkh3ipFNxvTwGYP/lPC61QWjyaT16SmL9cH2R4GWPCRrRuSltZF6N0DnkBEx
RDrP046mrWlNGQhv3ysKM3qo/sKVkR0VE+fcjvmEwqRCx9Uqh12/EuT8rafr5+yB
P6rjy7Wwf+jRsNHzIWOjGrwavxhuNX97S6uTwtxu3QnokvbdAM2/NHV/saAJuux4
r0DH6MqNf5zuPSc/hWhdwjDmrHxJ5I5YjAst/D/EE+WduaKLANxWK0XW/IdRh0tr
M5S4s4TcF4suohL1xlWvDFCEjweiThD6VtbiqM+epzVAoLycHAt9yZEQfT9EXP2j
GsXHEUBbyWcilj6X00MhGF1bkVJ+xWL/Uo8WgkSVjzcc+EAWE2rAUsa/f+/XxtF7
9DUf9KS6WJdrhZKkpS46Qv1ZWpiWXfAxx1SNd4HfJUZvtrmmYZZkrhwIVx+Y+Yxn
iu6h/Jj+NUjkPoFJz3d1ATnB7XnUbtZNLbcQasHtBjnw/6ZuhA9k+kUzeHNAGbvN
C1eKnaJ0h2v6XTAdlo0IZKqzb9yIcq92bjX8iwrcDdCOudH6G5Jv2ppTDJYNiwGc
mAR+OKi3U669qTMNnfcWpZ1Nony2DWDmZWrUrO1hs13Zcuj2uRWmGxnGFWKYiLqV
VrKmVQrnK3nHULG5IZ0axfidMuVvVKsgsesPqaxMI7MO7ysypaCrGCtVygta7sRP
H80gugMI4WX8j+bVcTxWn1PUSvVL3qmRj6JHzDqNrOgXOdJrxyEv3dEzx1Yocia2
XNyrSB+VOsKqB9C7gA8bQOpqaDckbsZwlfo/nXmD77AFBrKpSxZpZY+B8z4SVGBd
RVZlFP0AWMe7YQLh2k77mhbW5AmWVDdtIwx0NHtFcZhknQtUPt/CZGtp6Bv4h1vv
BjlxCUcnBFhK+ArqVGf5D+urqMStJVcqL8CJkhGYM26smHF20N3Urp1drK3OGRXn
KxTMLhmhMkH8dJhZESQGGqNR8QY6z5HDxKlXzwPclYYl9O7mQehmXaNzOspF/HGm
0aYSQ8phj+4ucmGPjTZOGg1wbKrbgupzwhcV8uEMGjEBduWs77qS7NxB7IZs0E4G
L5DpiDZH8IXhlruxZjoQymz5DKTG9dGJ+Ab1ZobyGk5Da1T3SQlhOaoNp0yHib40
GeAtJ3JBqPTT0fDLX0JmPFor+2AAqElxLkTHcjMcDmBNh6Ci//KE1WtlWFrPDyFt
CW9mGxiAU49L1J8CJaV1PimwaVozt/iYpC1kHRMPkdW6a0dpMEMYBIi7MbYW0kAD
lVr2NhF8DAIWX0XmiqfSpPH1AfTGqoXPdQ33Za1uynZgh4qN644YmYErYwefiWgc
cyXWShEayyUnlGSYAiSP94fB7e9p74wp4dk1KBiA+cdnC935ALjy+u2EohYMu0wJ
s0XSx+VtgZYro6kwCX/wx+/od1gekN8KRgNbLBRR4RF3eBlbwyeRUtR93P40FZjM
11+wFYWaKD0/JVNbYsVvmIIZ2sPqDmNowX/I5h8e/nGuelcqjuuNTRVL42rfvHBA
P72aMH3fRczOmLwvKsq8t7r8NM4RBskmgzo1QcshdxLfOrUyXZysllFRHh0Bwl2s
QOm1mQdGiUKpbCiZlvLeXRlf6O/kr95iHNcL52YnaTsakpMKzk6NM7GARltdxF8G
KH3OtSTFV8RfoNeZS5fGk8jn+C1tHaOXgSK8fn9gLZHdo1RFGQ0YakuHJDl1FS9l
gUZPLDzD6NaNV6z7DXfwI9zg80MS1bQ+D1OL0JWvpg80tLUdq0PunkPHt7LBl6N+
GE8kOv/m1f+dE+4UxPPVySB07+ZMh7gpL1vKDblF6pOcFC3Zt4Mw7b1enDAyNmiE
52nvKf/HcByfXNcWs1U//u75HEqRQ7mYCYmUR2M4t9hFz7ix/+Z8w5LA4Dc3IMgq
dQIIRHuVgcFFPRQHJ2qa6U+G8/VXwegFLJ+o0GhrbsVluba+f0bb1U3YE8Uj3aas
gGnkHC+vFitluqo18ZG0NO17VgQey3miFYqAF7HebDW+1wVflK68Gm0+cuPlqssl
v6vOyUselw6YbaDlfh4TPdSS390Icw00936dBixEN9/t9bp6cNKpp8cL/L+wfuzG
YAP5AFhQr0PgccFJD4wt2fpgkwdfCl2K//KIhqf/VckPYe4L3nFiYZBShYUXiCgn
MT37U9FAYE4qm0AZqy4ulW5CureOxWxR/cpeIZ5ignyiqllqGhDUU9Pm99L14Y1i
F+ZG2K1TqOIf0iG1Rj4HxgwkZYD767KO1bXsa4fRyddlz7tJtHgNPow/aIYs1j6u
VGbL/ZUuYFXys7tvcy/IVEuX0Z+/EtB/Wr1qqA8fpfNZCwbFNh3+CB0LvxVJ9X2l
ZKB3Mq7L9oI3VGHwKh4Hb4uNfQ4Wh76Cbduu2vpP68IN/t/6bGs+gWqmj4+NLZHJ
YUN5e7Cd+U/in46yffXw6Q==
//pragma protect end_data_block
//pragma protect digest_block
VyZl2SvRR8YkIJogBJkNZxB+Oxo=
//pragma protect end_digest_block
//pragma protect end_protected
