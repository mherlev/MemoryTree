// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:53 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
cdCieFZx36j6xiX5UeSx4NMpIoTMPpNaom9mt37PFy+qVxMcbD3nZNCzTXu2MapF
sRMzWcj5JB2RHT5ql24P5P8gzVtJcJdWjMpeFYmsyJMrJUAxDOMeV3Bisj9sQzIY
lY4feoGTrkqSoABvJwSs2sG3PZB0QrA9QlyngD77tB4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 31152)
g6E5+iBKJttgVHjUeZnYH9PCNW8rlv45ST/oG8UC71yZyqU2R2DHE4xsNCwZMisY
liCJwF5iJvxAN+q+lN+Xv93O9Yd+LuZwKqN/Ya5tIStXojU70Kw+B3Iz/BNLWhus
uejhvJUjlHBtWXh3eVxiKetRxWXN8jOWDD1P08zy/je5UQ74JfXoTrTnfQHUsgms
PpNBMk+1kr7Ll7/o6pDvsfXsICoQ0SNKoMEh2fL3BIfejo2Kwh0NJZCyBqJL+YRJ
z1Bwz3pRPhJLEfNN7eBiaAi/TXUn04K+XF9EA9yiyQ2VMv9HuMLPT5vUiFb52bmE
iOZ9UK8cnBp52rdP3ABRXyKQ5aU9j7GW57dhLnVI0gnE0whiCc6rSSc9l07StO8s
yvDV3hZNZGU4z2NO449CHe+NgyRJhkT4azrK5mDSn6mR+nJfcbwFDGqXxpWd/Qli
C1mvxCm0BeJSeyP/Uu/J2jtI6ykDEy3SeoHUsdw0eWuz4JspSTegSM1EsKWCUhA+
ee7o+gl3uSuEUPtVYyOaW0qAiIsd+5FxRHr3hZBaH31uWgpJwk5TlB/7RDbA/Cz9
Jk/x/664pTtE6OHQyMMrBrARxZmJv2U9LFW9aJz9UFYEgr5E22P8LCgpCsuT6cRT
rJsxt4HG6nyH9rH5ESffG2LGxstqP+w3PLeDzDzvc+MsDGUgUVQ4Omao2pqoJjRa
jHDA/qagxbrWwbmeoFMFVuTs4O5FJPxwYPFTVGxdx1rgoNLGt8Lo6TmSffL64fE8
A/yVY1ugdwZlwj4Rfdym9VPyig5D3FaFMX5Z0uyzuji5+crZLj9eNplJqeFzUdJi
8C3raXsAI9C5K7ctsk5wjfCl8iKgY+vtnEFh/zsUpjAL3M3Dx2z8EsiufJzjhjwP
xKM6hzBV5l6Nk5apqLrC26g3eaF6ToQtDPMUSbJ5bz3YEBKj2S0Lh6INoeQ16Ylh
IbUleYiS06L30aoBNQcmFtsk6ht7ExomtZwUysf78bLEsXgZOVwkarmuGEIc5/Mn
3Hdlk1Pv60q7TsfkRkhy2u8eJvGHRMD5hjBhy5kBbnbYf72nLITByjO1jcAe/s3C
IC89/M2dCNQh6/tMzAiC2UJelVRBP2yESNidnKiJJj3hkzGTcAKVGpsObhqsoHF2
QSsx9DPc7O/RgClRgPCWq3zM3IXaUWTUuLfOGxHsJ0hA7KVppVX60cN1EqJXf53g
8wghrPu4C0aN8h1haOquESla/NrHXOtV+68CBK90vqasD/sz3PpjWlz4Xupb14kr
jV7u1e3gRbcPvGWKLqFsbnFWCVydzMgpGzLIRdldhDZk2R/hwYalxmFgUBrc05Zj
iZjm2nwgB1v+TRtgst9jLfHgSJJsvhZqmlFGDyMGgLbIY8VSlHR0N0vUMcutOaWD
RfbZ996J2PbcszVuQPshXFXSN6/HgDdUxGY87c1L6wdST3kiiekFASuJ0FdBRWAX
MX9VU8dpxpVGN+bluYmQCEk6Ng10SdpVTu6HQ9NNDYw05Z71YAvLoBilWXfgVb1P
jPItlO7O0++bGL3JFHMwWe33FmWtc1wrejIjoCsXWzE0rlmLYq+/hFDUn+TatSZr
dEqEIDhGUG0HTBeMGXWrT4O0xGHB8FApiOEylQnCPEZU20eavAoma11oaN8uZtyY
ufEWp+HSTwlN8ycwkcYH6IcVwxurC6LOD09I7UhbsL/LYXBhLACzRYlXIL1Zkzto
L3SM6ZWkVmcezJ5/qShCQTrhI7Ry7BaZiuQmyHxoMXUUor8B9PR9BAdaDAwOJnhu
2pC2JuL/t3DaeWTdHl4KeSZ+5OYItN+iqBjNM0jRadQ+JfW0BfFHGXMpqsxEdpTP
k1+gBZuuyLvhz83DInfHXtI5kgTYD46lID1Y4F4W1ifHVvbVIY5K1MqR08MPh2/Z
QVUzzMe7WfEg8doBjW5rVvkj7r+Nl6hJ2HlJeNID1tHIuuxJLcGuQwOTa8zkiU3Q
V0sRPyI4yJVCXpSr4f+Pmkj2DNpgD+MrOEX8klG4nu9D3uk/OBOvDqlGv5PMzFgy
8WWDXqMwV1/hRhaB3QEKeAcdjjXl8lirxjTocyU8NcLqrUh5GY9WEQJTapBwfiFw
zV2mOjz6PE6bGG7T0icE1XG4Hrq0bJjA+vRdG00ueGZBSFxn2NCaPFCUfbYsqvIX
uzj4TEhK3PXnnlvCZ/EV5rLR3O0hC5Xl4Jf/C24VwIhzEzghhPepuPwzVm/BscjJ
mVsP3XW3uZekUrlj6w1c/l50e6X3mRN1LSDug07Azqt2v5ETKRhAtBg+qjtpWT1Q
c22fcIPGyvxzvmjEyt+QWJeWIHwOa0lTPdNZUqk23USDjwZlj1j073m48EIkqWOT
9hbyp7H9ESc6Wov9TuChRf5rUlqxsKd36WuHUI+JC6EMA9J6kmsrMO/ANN113hsE
UYLB0LK5tByOYg95ACULMwEML0e+EiDp9IHaFxqREXP7IjaDKqOCZ48H4DvqLnK6
zycdNK4U8vQLLWxKQTjL0hxTVIgfyXj/pTJYWx/5vqNLeHry7X2HrPUItrYgStZP
mglU/L6IE9PIjwWyxJGiDtPQ/9Zhw95AgXZh2klj8ZMbkHcACz3QxjATksSzyhxg
MOvsyUs9ssa5i4NzODwmsowfdfG2Dp/SjnT9U+dYRgyZbDZn7XVgyLjYDSpdv8ho
KA5DSwgkJAp8+uVGaFpCdY4j8vFwrRzrMDLdE0g7pUig7rS/kxWe81CMk0nBya4P
B2nPI2i4jdok4KHr06hyYqbk8Zfw6qD3ZVMQMoIKxSF6udIMtcwCiKaLeXO0H18s
y6fBoXAS6YYq4ptka8ZQv5wJcaDUDTjT+jCdvtPMj65UffUB0oAg5ONfz9g3VEpA
VFt/oZODsiZ5l6jMA9WgyZminmrvlp9lgrAchjGD+8OiyI0vbfxNvEDFcIeA32hJ
O0OYSp3VEsaFZKTqtjeOuQvVOiJ0JQt8TPNYeyAH9hdKPE+S9TsXpmWh3y+C+mhs
EPyBNMF1DvIj38hB/lflNSXbJUMc4s8pZoHqquyYVIS4JCYAmv4fQG6ObHxpfmRZ
B63Af5MZwJOF1zt5kuudr7QJuKUD9ubItce5WclDjvFPJepYY7wWwi3LecVC64EB
p8zE1mcRNQNFB8/m4zP8fsJSqE7qCtHEKoWy9osyShTqOzc5lKAHNARWjaNvBkJ7
rud754yQhhlW6x89jpMVXdmzIVLQh1uLda2U8XVpgk7s47UTDjVmQCGPJ8vQUn3i
Tl+OUQS1A8PKfnZZ17VVBY3X5qf9E/6Ryx97y82ecxa77kdeGjcdE0l4YHJn9SAm
ECX1f9miEZtzC4AtDIXZ1cL+IHMzQA8yOMPHGvp2/Rth2WKLRF5YpUBOe07TcydJ
YVknWAQsrWq49FdU1BGn0iSAdpDbYOaU+FupROBCpI9Y57qOAy4yYX+fsBCvD+pF
vUqqcHVJfQELsjCRIOq12Nvc75pyM805GOMFcWrcG2jXqsXe7qH2PHOxl27ZYBqV
xvhRSXSGPhbsjIUjOfPIVK8Eq5RqyviWjzZrAa4oIs1yQO1Hxe4k+Kxyl1BCu3kx
1dVOYPJD9NcLwuYGJiLkFeGar1o9k20+azaZpjFgvHBjGFymAFldIONT5R6XBwfA
n5vj59CvrTwgufb80uSQA6hPD9OmH7yVgjJkKIapX6dAIb77yoLbTzlGzzDBuXkr
pqE0G5RQ3J8S/TGK3hun0YdiS2X/66LsYhJgEw8OGHYYIEkbasWRjTU+rXcTR+52
dIoy6ZtZJ7j7AurlHIw5kHBUuPBdX1qqDGzcV7pZXtdOusGmLR2E4JQ28gaZ5pms
L1mwmVA3isznNzQe56ohJu1O/BDjn++bfzwZeoLgFHSgk4k7+pfAueaiEtUdLyei
tRaIjNHcUFF4zH2wE3kS6mEJ3ROfV03Cr6TAN3Ol4m1R9rT1QQlVSP81KiVNZmk5
giSmwSND5KvDV7fhSzI/IS0tjMn51dQYvB1/RqOtjiAGLcRPMgWQSw/1M2wsS9ao
Xb0qMbsNViAU9bxfIu62iWs5B0t1iCN/NagLhlyzGlC38WnPgdggiOZfL4/anEUf
ADQ1srmbFokuBWI5Tj7dM0m5LhD4oE7akrnGpw9aI3aTROhMIvpdmm0qYHvE8+oe
wWlQ1Pc+4sesFh0YeidC8j4KfXd1yPqwIilJcJ9OIfGI0hyOtcFOCBeNYupUD5FZ
VXHs+AMDWsEa0nbVgpyl5mdlcMvmJqAm+fj6RuFdCP76lucKgKW6gk4IJSV6f0Rd
C4gQpKigK3oeEEc3/30LnEjzUp1GvE4nWwVMPSXiMEipZXehat/WrW/YEGNvkjcc
hDtkuMMe2b9ufuF06RyVxvQ9WjZUJ/75CafsW0QmEzn/al8MlqwQWhDzxdfwjToX
hp1DDB8mjKelnkhBHxXWnd627qQM+XZMlqjpsc0AVuoihvt6GXYB7UDzS+wjoVrP
7vjEjhXgQP/A5W44hzBIcMcB0Bc37IGuppmkSDNnmTMVKwttSqTDcvtZe4QTZmqS
Qde1HozKkpLx0DQnqLA/50gJTBud5O3QgcdYBvYS2Yb9yXcKQX0luF6E6kEJpxfU
AgeD9Jrei60AKYztbAnTcAul/nsYLgvYbyQoTseKEf2niH/n510d14sVrxGtlAU6
z/WHNyRA5zsFeG9OOJjycL1JtRwaW5rDL5LiogXelST0/Jp9bjhB7AK4nW9oXy6s
tqvjLz3slZ2DVjG6B0psZqwx/xBMuUB9BKmWBO0znrTWjfn1GF4cKoPTgMmD4D8A
ogufYu/WsfzD/C2h6rgWfzg3ngJ5LugswH+RR6MRH29GbZ0THbZ0gwrcajNVuEbE
+HYJAxicqqYAMwOIC/Q+M7WmlzgBAa1pkhpUKbNfZ61Vu4vHGyUmFuI8UjbeHckz
RV29o6bkYB2qpcB0vKb3b5eEpD0prtrmkmfdlbCWFnF2GGtBoht0DdnusLaZ0Ewf
d8W1y2lXv3jvtAnaBUBi4Y3zCUguSlaEuo75zV1ly4TLl9Vedh8JEljxeiPh7RqD
QK5b90msr9tGeaVzOknyVpeuz9ASpDUtsg1agQiKJIMtggryY9aM+AUhO2LcJFhu
dc8MP2SxTWuEw3mSOUDiz3PoHDGx4nAfAMbSFMDW+zNPqFu3fWZDsxIsYJYtiToW
g1ymmxEPVs3bgGbc/Bdk4IJkB+jMJyLF76eUH/TBDv3xhWm/6ntQf6vs61bGECeG
0vwUgIHyIpNmZdmnMkv4lBaUpJu55v24y2GQk4Dg958WpCnH/SSi7MOHyA7CoteG
mDuAR46RIshHMr/U+8Y8+gCW+g9kpFc/7QmZhSwKx2qg/nAZiBSe+DBYNIsQAYk7
dPMRGwFLDZkIGI1OECc6jAANd1koLknaFeElVTPKcXfC4WJHWuV+GTGYBJoAE2QF
y5+nkuqjen4vJFhCsTSPY+RsJ14kMltFBgimkg/5L++klrLWgqVbAHHPmCpjBdVE
5KyzFDiYKdSJClv4f6K+audbRs+CnZGViuEnX4sbKprBQ3fgt9+9LJl/tquI4c53
IF4yIQiBoodVn5xu6NP2nnlgQ/rye4cwxs+oAAjnzlputGtdl9a+hV4i8bV1jktU
ucdL/l+aiabttzmdHNstsWsD7PNJ/mFxNcteSovVTjjL6KwkL1SxowAo1Q9drawj
UvbkQ9ABnR93FXg+s5E9NkxpSr766xMJ7c8RlVh4ONNAecm9xyZm9pLHD4TqeGG7
3K+1wXjH2O6OTn/eu31f7i0JqEdguU4auMCz64pVlj16JaDxUQ4shF17dkZenmtb
FQrW66h4LVKaqiCn/mdmg5/4TO0914A3Ok2DIwhnoptIz8fwdDAlBo4FkueSnh8G
t3FqV9/Sc/jnYnN9xVCY3SPUoGqQXJXqAiBdfT0AhQMOkj+mrzduvM5pDeTj9qiM
Iz6gDc3QgVcF7UduEeCpJyJg5/5gGEeYRfVxkP2Y5CF4FAcPBotGOKpTWfvZ2LSt
q3EcXkoZuEp7Dz60SdaNWOtw5yLlHnr2kX+znXFQEemEMZNLYrxIRni401qYNUCr
n0btALdVTwgsv18Ramki73jGfTGzyReGCAXtd4roLpRTIbjPXaxLHctgzB59nEoO
FvXqIaQ79GMD1m0j4/Sl4XgqsZGo13j47sdb3oQ6T1ertoXb2T94A4jYCsS9YubV
ATmiNfDb1b7y1W2XEDLoCtENFSSOzo1RPMO8u8IJYVyrWteigBIYzYHpVBjkg/5k
/vtVUxDDcFDiS9os6XWuUZ3DIRe1RKA+DFYuwKCsD743LvZZ39IrQo/We1pFAmaV
F0wOT8aX7b8Ko4xPWiEjK8t9QYlbrahVMOkMst+b8nQMaQ9QNieRB7rNhLwONn4R
OkwSqKsBQlBJ7ncQan9HNBly54MDexjDr5FY3dtnPlD76MOoO28DtdIlw2QUKP2y
XZ8iFkDtCAsRIRQIQHq7tTowUxv3eMQ1R6N8RGIDKzMabIDuTM33M6HWfe6kBKVl
xF3RRraVZyjARAhA7Rd4UcAwxSI4IdQuO6G6wFSbMQwHJ8pcfqivGrbMNzXYxdVZ
M+DYNX8eXO66ldEKHXcqeb5M3W51cmjWJcU7siyzt84DnT5xUb4L4w6EIOeV1OOm
2lY0ItzHEvTqRAt7huvsFYsjvnDmIsTSRZVpkLy25ow5aPCK4CK2Fe2/armCbewa
pTrGFposOWpe5p7HiuIpjaeZIt1hEk4XAv/CeCCibfnZU2cR+6WUZhStbgcfGGp3
87yGykLbOJwzcC5bjE57rXdOWFyIGNeFHgbEti2rNDRlWA6NlDEaJQduxi/GP3Vf
6UvGuf07dutDmdkeGtA92SHjdrap8ecO20L2srD9aBhEflXDlFRrdlQtZaFcwMEk
jEsADrBn4JII0MovpQnVBPIVgLqsgeJBD7UJupeD7sQrhE+NkCDzXervMtoIo8DM
FTZfjxmtnn7ptgkKw4rOmdH2mbGL6WQOYgSo+mRJQR/AJEiDm0bM1XkXawnghG5t
uHuNf8ba4uifjuXWDSKxvKt2ytAgiZM5yua8C7+RlunYu69McUAqTKh3FZcliJPu
ovnClS2+a+tNrIJ3juRdZoQmQ5kWCLYRjTAU5gcuGjhxOujx1OnVhRLvg2gkn3Y5
aod1uVPV729Kk/aJeiGccwkViLC8K3Vsz7kVUFGvzCci8OWPUsPf85OWddvX7FaA
ydt+8DGgftdlqi+Vr2RhAmp7hDn4NiddYwmlu/2IHg8iluLKw4mdC+85MP6wa2Uu
NdmdUI1/Md54ICVhiFqO+vmBLTLHM/5RqX2HDEitZR+g5Vqgq2FmOefdxF2053rJ
k3iodPTpwBJKehF6r6bLG4qcHpldpNUanPdAKFZ5zvndFkzb3tVFVJAc1bKARgFs
P9RxAzvsRoEauwdRGuNQsM/f0mUc2p9OysGFcIlMh91j6eweZAydhJNZqRjucM4S
woVhvMpeR7Qph5Erg64a8y5THv+74ZCu+COle7T3aoZVqJcU70FvJ+hnAlDzWCu0
fbDON/lYPGfu6pWvC2/Qm6314gAmFKaJZRs7Yp8nORv/9j3bK5BWY7vg49LOqdOc
7pvVEuXVV62Qpz9P7P5QdKfUi9SnU7Xf9Eb088kkCntM72Y30jwHaNsyVA5klvWK
inwiUXno4OboGZ9wm2Eg6WrT3JCgi3vE38rRM5Rq9Fhb4AjYNo7MCno+HrUuLDIr
rH2cIpTshpn2p8AlAvw1OZalDIf9QiKPV9FQJqfUVsljXHzG8mYcyKaHJ3eVG/A4
RVNAuBg0KEOtGh5Wu1IY59vBOagSd8bHc2xxV7Zbs6g4yhBkQRfhKjQ36/OflGJV
yv+1NgOAauaaOcwCoIPWP3YynXpRVSm6laBwM2N4S5cKBVcOi/ofZs9R9HOQPLyV
MMHhX5gT5WQsVGeu6IwF1ENxnV1d9mlDanRe9lwswnmKgupV5OrUpoZMI5q77KtQ
zsa3X2OzdLXAuLIriU/TG2zkcdnvyu/ho4VcDRyYSKerlf2o0KIcUZiE+zspxb94
aBh7G3MVTl0N0YbyPY2zruchtADGWuRDKoHx32v4rP8amu5s1j6u4yQcLDEKKx1G
x0pwVCO1euByxVgU3wJUB0p5TLwdNshGWc9n/1rkceN9lgJj+wiWMyDI+K9TrA0D
ESxjMThq8dBAi+1XF+RWWYHI2SiG/CCx4O6ih80R8ajY5qEIaIhfI2v7+XbGECS8
jLhvVZWPXrORO3JWOUPVxPO1H4RUy7eZsU/dOFSBjBYZXusupHxPY7qX6oHf440X
2DIfC2pBrl/6rKrSNSfMGOVHSP9uWjtCpkd6zGlEZ86LGO8gnYnTsCJohVh77V/6
EACZx+45IQR0hpw4aF6NmZ2k94xExP8D7Lpe82P3O0m1ENc4g71Gn6mWnr5xousq
1C8Gd2/XvN51sIO3t07S0l1Epn4HSnQeDOvLavAFVLWeYEg7C8I94Ycm6uLHYU7+
rbfOeqg2YSGdSnTxG67fITDVKDuSjNKox3QasJZegmZojP5vfNOD9VvsYdaYJ1sL
JII5rJilacC5GGwMOtyeDnoKXnJd0mFU8KNH8qPT2INYWpagsnlN+yIE2k7ojpOy
2mNsrEAlCzT9ddGkbt7fc111HpSPCxkgrKEn3AZVkSpxYLG53LcUk/AhiZGBPa6r
UhYy1yt0Kv41LoX2+Gfl7ZgbsK4ItiOAAeo2DmT4JMVTyhYomdKc/ciKdytCsecV
hccCV3NVhlQ21x49p734W8HyZVz2QpKl8Ed1hb5cYQE8pgdZ+MSpkASKU7aHzG5b
VLF28FX46TD6R1WWjAS0c35nZG4SzDUAYSlN8Rdg9c8pZn0+7KXvGJCK49qvYP24
AmG/7sBLHvYoJdoMD5S2hL41eqqBDdwNB4lhwHFifPnIzUyAE27O/DrTJSQlWm9y
TuKLfTGG6MMw9H4Z6aJm+H6FSNyrgSZDL7MyYHPxSYOunRkQ+J0q5aX69uxOQCMc
X6fdDKYm8uuPWxI1uFnAOmPd9V4FjOPQhikqpZFFbOwjePz90z9YKYmzTMmBhO0Z
TJjoDxwfbVVYT9H2Ju7cbuYvfhVwy/DCIjyyC5ZCv//MWn42VDmqXPzZXrcrILDI
7TO85KnUp8LtcW2eTJSpeRNKUysm1Lax0gOfQDjxknXUe8g6n9LPjny5ITE9Q6jq
h9l1VQd6yfpW+6zAAc9x0HkHl/3Oahur7SpDhHFRXgKoFpQn1nUIhYaenE0Sdibn
LWi4SoNB46qBmGWYex+C4Zc7asGPhVPqvYRQwejiiET335iwllrO+9gmAhgmQ4mU
p2TD76nimFu2uY6f7wNTlKjvW1A3gG0rt4B3bXstAPtLSBMX6vkZePwymATOQ9eP
epB7jZs9TVQgGkTX7xKCyhPZyEQOxX3zn6YEtLgsMwyjAn+6oCwdFVg3yvcsl1pY
9NJu+ewmKVjEQZhMKeiyqviuAhOJDkFYgI2knv2bvpxdHUpr88wHYAVAVd4efOdD
GAeKENOl2+Phadu2PheAPIZmKalx5kH3lwNsVfZ6nO7YQUu9DdLp8lGojjWuTIK8
FPtNpeVFqtM0mW6ktaoR7zxEWkm59xd6X9fgqSsCAb8CpNAZfhIg1t1kEpjFHGhj
Uqp1EoFk/h27dtunwb95PAJzzEHdpsiOEd36KXCLSNYOdQbPMrEEevwpGZBVfv36
wY+qyIsOcQxEAeGOoXTxhu9gqpkpUdbQ3xApQImsYiNnNfzrRFlJzxYhbDXLpVd9
wl8iAmWqyTeXDyl/qi1uT3qIMd8LWNfdjH35HQuuvrSVeXpkjLslVdPeHPWNZ4TC
F1We3vdXojPvz4vlYmh5WiitFsnrr3QnaD6acHvAhUCMqhdHX1Oe9wLYQvV6e1nV
AKkOiCAICpK9tTroPpy3EFLT+ocptOXeZZr4t8TjedfH1+cSldVeMbUtxjlKKpNR
AqQeUumMtrz3AwlrG0aMALSe5Jn87NokMsoWvJnYs1SLdRHxJFCO0ZloJ/22LJur
ana7CYwHq8d1AMUeweCE/8dnnlMbaal8ZaFKVF/1zin7d9ax/OT/rWW2P/raD9rW
XF1dRpP67wdBfLjjh+Q3A6SGkR+NzvP7TjL0pHic9bMRb0gfW/f0Eh4vbg6bD1oz
dPPZfsiJSYv5pJIYU6eU15WshakF9zYropE4t60ooakir6r0NInTrMiVZyaHv9Ig
KzyZnrH1jJtYhOD2nnVmcqwHI5I7QBwtjUU3OlQGyt9h4Ie5pc1jpmwjCRzS10ks
6Oi0kTtyEcXbPbyxPwzADI+mvY6SITrpCI79+zlajGUUxY+DGBrysJDMX8FSoAcW
pX0QvCvXy6sixu3GCbBYw0P+3Onz1AuyNjO/xqJ4cFdWTPOczGJr9UFmX6mQivUD
l33PxHVpEwBrHla+m0Kd+b2QNDFEarvusdjP1HacPd9Hwr888PCTplTsG8MfTd8m
ydWj+81PmbUZ4r+d09mNAsiDo7Yku8FIMjtA8zHou35R3zNjcCKLuUF+Yp2qaP/X
Lwu34JBPjqtk3NhgNP/r6Nt0+Rxda32gyDe1qxF+DRQAlk8YjOlg/zCfPZQiRe6R
CaTbTAHUG5M7im8ZxeJxvQIQeDKMxDPuicbqnWrxfH0gkXol8XG2Qgoy9dpi9nbB
E7q9q1SHFoEvPdpANeOHKFX+b0QhCt1q72Oeb4OOiYRwoE0r2sbQPgh2+jIMXxWc
5aMxhHbn1/QmM67XjOV2aDarqzohJ94cK2YYbMIfDdpxF02RfxDLbqB6gxOP7OkC
2u2bXr5HcgP+mDZNteWkp13836wElkGDK2lcjBxkBiTF66VWozbEt3LrAcMqGwKE
Mlukflj+Im781RD0mc8BbCsMcP639EoOT7xxYLcHHP81OnmBuiHOnF6FCCxdIINP
TMgELIRnvIwMkPZm+EooqAatncHS/DgQAxkU+PZX5Dc9WtKg336InKjoYsZG2QrW
2OkW+TnK1CmSnjzWuU/tbOGCWVTpoGjal+8+u9ijLPDeJz367pleek6KlNf25BeY
VIl/BpdRm4O1PkPxBsG2h0orLgL9kovBA4Ikpdw1Oo1KtgOar0U+8jqCzGpjxK9n
9HGAb5ufdCQFTg4r9hqrrElPyReV8UuCkcESpHKbaY2tZAzoXRo/hvnRxmbMa4VD
39LAAYT0YiHMfWpWU+Mvh6AL8xjeeSP0kVGTtyCu26sfm1mxG55agIMgXxywpQyW
C/gW3aOwdlf/BwaLez8qbZXrms6DDBZIFW67NIwcWyWBVNZxGwTGvf+kmqE06eiC
1+EduoFkvz1oo5jML+aeDCMKx2eUgU5MEmaaxZWG72+JrmmNxn2rchnuKh5uGkr/
KUk1GBpzWP6Iz/FeRLigJr4LB5YMWik9fBoK0NBdDXCgc6T1CfdlqjWCPuwCj6IX
nWZMQfNJcg+KcjyM3kgkAXkWfGFEWeuqrnrXDlZp1tFpXlizAHha2rBgFZibRhDD
UXFYy2/QSACCPUcNU5wkLjtYZLMRjhejhwaRrqyuc1w8vcQZcPOmPosgIXqsOQCS
Dm1CNNDNFDYxhBgGOsWoSgqSt4PT0ka2hkDpGFFPwRnAaqvsDNDo/ftJLqAWaRVU
d1SmbH12Vyjbyq2iYmrM8jvUggVXa7bdM/uTLI2g2wm/fEolUWRK6sMRbSPtEs22
YgWY+y8duzcK0If3WbZm346Am/ikQ1WGObyZW1QmPYBVZZSU+R9Q+TLyPxC7kfy3
hfn8rQBPDNgiQ2Tuz8Z2RXyCf7ns60E6vELps5qjHhtffUkZiFYcMlYjCHVCL/4t
I64AR4IrUDSxQg7TluS7CT5JZL3xmnyA06Zh7RW8IRqg2eYtciZgsdEpE8jKir+R
1fFh9kjj1GZj+1wejyYCkJv8yotKAa8TxuzCoaIbbn07nSKR/SjAV7t5Ey4nDiwL
MWODRVXu63J44MFksaKW+XWx09UrAz3ZJC+7H6BNTNeyyyuqO1T8/fk10/OXBfTM
l6AiXY066+SFenRwQjmM/XNX6E2hOSfc9zT4qACeadPaRqEFRUT2MhhIxRLdCaW+
/wqvyeomaZap0tmGGAmksH7B/Hlwj3gHzK3zFo1oFLwKGaeLSvrv/ZEfdekzhH/m
wANVyNeYHCW+Wp+o8hOq7ybUh9WihdX9XyN/iKnXBj7QSoe7qzfMZt5zobwwZbTQ
H1nhrWkW59RQSyD9AvBiBaqAdfGDSvgoAhvW/eNYubcXmJpbjI/RbwJdcS8MWuLl
KacSw7+Sr4aP8TrYjoj73sTa/41wgqXoSFGUpJ3t3gTJYSs+bs0kq6yzzuA8ZgN9
piGJ8IWv5L8O0rq7KLK7RL7ENyJjbCWJb7y383II8zQwbf0H73i2R/uJ89ZkYub2
rEEOAajxaHtr7iyCiMaKMgoeup3ZjdzBLUxtzHQh0XQ+0qzpfpHlLeELfMHYLCSL
34N73OOesMvXhGwRee8v5ZLMs3OBKqRIXDSP21pj87QdSZ+1Ony9g4kB4mGXRo//
Aj5tECfAD7KL+Mn6+cDkDBXUhqOmOyrFWkNyx0EcXRJFue8g361/VRm+xc5qOfb6
+YEg/0NQo0d+gkDmBW7HBsDo8RzDNZ5siWRvb6GBNTl0oa1SDF9DV5XmUZACWgzB
gxpmEBvxUIsSLCqDiOMqIC7a2neKZ987EcFtJ7vzKGhvSa47oNAX4CrgrQwor99M
byux6ed5Xvq1V4i3jiXOBQoGptWeoSN1mefYJh1bDpgft84BunUgoAwwxYQ5XL/F
4rHsPtU4UZpUaqyvNHTPDdcfYK16RlFOUH1layMktBhlCwQIV3Rr4Ds+vYM9lCE5
xjB3Tg0rcz1SEcxqqfk9LXC3sg7S21Dyp5gQUKjhQhSqWUyHP7o+69ib7+oqJSAT
gDvuBUwymvOvet+KG5+8gHBCvLz8cNsiDOfGZtnMJLd0EGeiaEKW52OrIPGh4s2s
gAY3VNxesHbUMnzlNDqwt0G0hxOZgmhfcuzBrPOGADnzd2jUXs4gyheNe31o1VuM
ET3Xq2C1Ue4lu5txzp58iKNMXsH2T7Vkl96F/OckRJXjPYTnM7LruuLpi4Salv6F
JPJXrO4s4wTICGlGo3EgZC0k4YUZGrLHNd1xgJ4FV7EI1k2RaydZqbHn3JR6TdP4
HgU4UXjLkjBz/QlsVk1Bf8/cl2NVAdWjEqwfqvVUAd+2p4dljqou5ST/DNQ5yOXY
o3vlsW1niKuVRn1VY5ji+A99pK0JVDrm5Fx8qTlr3+HDMEe8tXHvqFxblGl9IbDp
lwcrmVTjr7Fa8DDJq2kzp6miqGBWMGM94iz+PDsIqrWxQmHnrKk5RUT/eHC+BLu0
oSek2T0ogMzhPIA55gLebE0dSu681mUjp8n084hWnCnaqP7uMS72rhQSR8QeXi+f
d2pHgQXjahDBdXNHPOvHqh+DtzzLMGyvviQrKw9RQLVMJfiTeQlB/rEUyLSpycP8
7HO12Yw907JANhKhGGIB+v2BQjWrKLf8a7YWC4Sh8Q9mpKutMzc7OpxNe+im5Qf8
LTPYfZ6t5hA68q9TtQK6jtfgGvKx/cI7E5xRzIsrYXFiwgfvab/0jKEu/UR98FWA
gLMAB1mEgvtXPA5VZAGUeB73uEZ7FOwF5CMGTQtG/ElIq5eVFyxw3ZQhV4ds2BGu
JIZjn4TZ2iCD7CnfLTZuUnu1JzdGxLQ2Z+CbLVUMUKljkecK1NJS+LEWLPHb8r4a
HI6fevvaJKjra9qThj97j85qNU69y32QKR91VAAEx2eAG5AyB4yY3W1etVFN4chr
5DVp/9OmpZdom/sOJJ3E1zP1SkxuW9Vd+VIywNQwQcVhQoxSxj1amPSoC5AF4NT4
wlJPwAoxS+p4xt2byWdDcTep8dJ8gSSO1ZiyujZ8ATosZUZDXIJQBKge6/kDygp7
5tQ57YL/12gN3G28ZC6FZRv5pWU4t2joPVJbdam1VQ7zGboQM7kVmLL+2qhaLoh3
icUWpV4jUyCEzrMdqoNfEnc224ppes1XS40gU0yPBON7o1IOLTp7n19tgr8C8qp2
I4goouQcEQGa7uh0moIaPnXpT+Nvy/rfrFVRbGdolP+zcj0fhmxBibP5Djvtpqju
ar1CjnFdpgZig2pR8YJHjpJBdynfYQ56Sc02zT9nD107aPUJyFd01wlocptjkkxC
0LK4QZmolbcevJsy85ZVjKNGXXl61wNHET+iy6kru+prLe0fJca17kURAx3GmaW9
ST7MsE6e//I010A+UR8DI/jzdgFcy+LH+pUyJhdhBEcoE4zlFJPg+oFBouKiooSn
1X7UL0g9kf2CLLgLBuD6ILCgZ7vmlz00PLjjWxUCpjJy28c3JT/drTWsl/PKbBEW
k1DnNXktMV/3Ssm1bhxf2AbZVbmR0KN0hRqRMdLPjwdLAVzlJE6+Y/yxZwzwoydm
v+hRQ4deI8Hg4L6KCRW5OdFPcSVDR9zpDiGYc89i4aO75O0e+POLunmWvRRcN+zm
w+w+cw56d9YXYVq6hcrDf74ZoswFQBiA3SwqND5WtVU97YeQV8cj1Nef8tgwmKOE
k1Sdrno0Z4bYIJj8OHpgQza7mwOjtfVbf/S5Q9j2IsOSIgVMqJS4XmZHiXQj2rEl
W1Jlq54dyKyS6C5okJE+Bap19qGMYUwprGR+y3LhjMYopMGsm+eU2Qx4x0kDvr15
SgZXoyxAfREUzFcj3yrxiMWpfawwk8XR0PCn4Qo92hXND62ZsS1hxPh6O+y5F/vQ
s122g26yQ0yzF/xD5uln1yTkokpDyE4V+5PQobn+BCXlFkA/Hc9mYG2wnf5ZT8WJ
SQVtGEWbb0MqZdcVNNVPUKNCwoOSyCfXSja/txMmJg43Fo9p7T549KPoaTeVTY9W
A+ch4WCVXqTWrqB23R1ZHdo5O+t46XIIkyq+9hTA8upDuxhN59k3+K6UC3jEoQ9l
UqEePppgKYtkwjpkn2d47OzRJ6mM3Kpn//YOEgJ0rjnydAty05Qm06EdIyGzF/d1
ltvekuDobK6NDMIGsiiRTd5WkH00/TX1DTrjlPnuJ1YQ0yhQABP0EOeLmf4Po8pK
xO+FCIpaRO8j3L3ne6mN+rQjb0e7RMxMEE7AJSZvsfapHvh6+yd+iTRr9W9eYW9g
g45F6t8XXW3FFV++6e8snJxgXsnbYK07E3I00cpaybCRr48Z/JY6zXkoaJyHkjGf
cgk3B+ZHyZQ+MtoCW8xDOdvORvOVoveukckYfXX8qr8Lo8pF+eNKRPu8feHq6vyi
ADXUmS9x2iTp8I+r9Vjxnk8sxS+9vRT7c0M6zYhwEFWpyHywAkczRH46zOGNVfy8
Vp0omWfQ3wKMmaTCAJrb4r9W4YcRDrAcLtGv6C08VwwejrTZirkDi9VR7AIMY8sS
+PXBODWAIdwc3u9Zake7kOTRI+ekOjGFUPgjmGrcH3tZndJShdKULYSHtqy4pwU+
sAaAFeIVaDRc3sn4LDv1C3cVbA3c15uo2CNHTv6EoXtj7+hiZegcTVfCgHNDYwfb
RoQXy7TmKWHIJcRwjb4EFBtnNN87REBT/YkV/9Iv4GtW2ndQNWm88LoP9U/fNZKI
S/n1/vJgk+MynTQxQpIWdfLxs9h22UGmdbJIgi26H2p2XP0cRR/yJreKqvrTOt0J
sZJNw4cnvjG8iz2GFygCWjxUG1cD9j7jCl2gsL08bZIDX+P18oTkH4eKK6+u/mWc
729XJQU5oWidvmh8Jv7bLRTnyx4FVYMUydOhyuqaaOnCaeM9CCVK8Z5x+WCf/v+h
t+I2VDXrahKyRXksS8AAmCiau2H4X9hFplviEeauDiUU/Q/66pQccusNtqmQ2/3/
LGZ+3e3V8DuWdxKUFnCXj2pQ0xUvzpGV1N0r8fJxAyIgMU2fE04UlvohdwxDyA6w
MKXH0y/sO2+6RIQva0ulwbCi7hSokdLjNG+HETagVlOIOZJnw+sWng7L0Lb+Q980
aQEU7ltpns3NDg7Qr+hbBVHEWMgdpK/LKIsBeZQ7c6P720goOSIDIDN0/yxqEGZD
5000ueXP3021fIlhVPPic1ItIKmCfaF4/IqPXlTCq43+hNAWM94aMv2fWwQcr3iy
do7nnVdCRzV8MFkJRLeIwQ3lsIqQHfmWMp073c2kokt7AhAXb0TSS6zKyuVyE4eq
MLyZE+XE8Z25SC7BBo9JSpIdthpd10u9/HxXmAVowo7VmCOvOmKkAATXGvcQru9s
iUdzhyrP3lZWCKoIY1RSs+QYRazuQEytZnU/ttqMejz7RXkUAEzi1fHV2+DDw1Ir
JkRKA7wwfkjTD38HuIyaKRHRNWSVnPrNj1owRRq0xKVpHv1q5npoOJPiCAywj+Zm
2PQnuVbn9R/5xEGv/NGzQUFys3xuMrGU4NyP7kMQY2VD1jDqGzU7230vEq+zZfQX
nJeV4CQ0H26dToXgDiFrGJpio5EKndby4zpm5Gc3SBCdjV9RFzDz3UO2WPxNrVZ5
OFE+kzlRvvGfBPMQJVbt3VOXUTTQT0bR8wRUm9KI6kmOpclJJigJKyJjB/3fwZsv
9hQ7UKBHQi7Lqv0cM35qBx2E6o9UyJtbDny3VWv2goCUIdNiYmSuvz5JZsZpSeKN
DTUFt1yOznZvB5YDDjobf6F0R7768v+sqDzplGUiAdVgfYccyFa1l+xJyv1WwbOj
1ZpzVd+Y4NFJG18DB3AISsejXrJquPNqwxEoTJ+zHA5lhoFI5k2TBPU2sepvZVXL
bWp2SBvs2lLrfn0Jnu52IzcB7PcmlMkQ3vNXj5n0H674o//zz8MgommeSxrfRJXm
5qyNhI4nP5WDgGRdq9koPVapG4F6qwFTD7J6tY1KmVz6ft+WGXf+6dSwvrA5Ic8i
LXw72wC0LH31ZTABX9E6zcOaLYCIHKlGVKwLaSnqpL+jhkxtC5sBOatOneE+XGon
7pyFaRHAaQgSFdx7y2QZuLLG8TWE+Rdi+EvkU1b3UShUYS7p/8q19r0pBpeVoWJg
Wkl4Y717Af4XhZIgvOkkDEyYz7zgbos0rGeQzL/jEhT61guediKkOdw0K5fl9Or0
oTDNO5HgN5au2zvmBU6aJFpog6McFL7cKgDGAr4cW0j6XcN6HESc95S0qdmnf3F6
bXji03S5Aay45qKAad2R9eJpJdlfYl4T7tVcGHcJ8DaWGs6sBvwAjS5XZjWpbbzh
y9oSgQrYU6cfHzJ/k7Q55N99qEQPDgkgfUbCxA5Ey67a+kCdW/jeMAv3gQbaKiil
avEbICnbOxyAdWgHfh5tTtCezXa0DNA93cW2RskXkmbbnzdRTzJiF2o6BSWpSiuk
3HXbdPLZz6WBuRRfgGZzKnQxqcuRwM3sYzyZq1rfGXhFBSXlQM4ld0txnHKvCUeP
aLPtWNu5W01eRZErt6+X8Ox/fXsdr1nzRv4cRYJ8bYHj/b/BBkMOib/u2jIoqP8y
7SItfY/KV3F1aLHHT3iLmFXBaDh+RwNGuFPU/P2d932lLujbtEL0BVG2aSlg41Gi
+u24NfNYNx+hM3mUCRQvR+XD/nXX86GQnUKFaZCJhfNyWFpM9n8DWZQxSVMPkXOH
AlYowVODOfyVXyKoEOTr3SHH8a3KNvJoR7J0YBamTWJ4nfqhgWAkqpnfa7vDKjrO
hjJkBb4INqg/A+SPvOTlZq2SrL4nYf8qWPRhmQ4cAEDF5a30AVw3juLR2C4t1F+O
eo63wdJ7qwFz8GOCn9f6Cr1Cd7IWm6jpNSSyhfOZvR2I522gk/W5Y7S62pmTY7GX
KRattVZVgC4RZZMskm0ksXpvc/ZFRuWgsDsCoVWalR1haA+FYKsxy4fYf69ztpGj
qkxHkdS3RJiHWpk4PnGRqu6APiZGInsrEBhE20Xczsmai/2OcqliJaBsQmo0e7Po
Hu1e1iTAZzMqbipcE0Ils4FTtdrrbUDiHrI6KR9sqFTOP9k6GyNuLUNtNIDCi+W5
4PrVshDCVLFnCYRkgjE2dIHQdiZx0X1zWC65LJGfmhFAi5KzYKBDMYr9IQpH4lKz
Qt/8OvH9JWTpFZjl7wfwun2qMVsz1yyMV8a5ZNI28jNKxW3yZKS+oPm7zc3IkRki
U5dtT0Hzy9mzLxwu+k7zNvOuSuvNkmmwpnGGy9smhWQgnhfGLl0T4+oW+0pxo4DY
nTo9Osk9tV3rWcTHmuP50H6GP42VG27oHywpOZyhLf60tjcovRpoxj+ecgxuw9xo
FMQJAzz1P1RugV5l0ik7YAkT1owaBbdqRGVQuV3jgD8EdZXnuyQhzriYcEZvk2p3
TiWsfGnzg8zgV8iUoNNyLCOh5fmxXn5a96Z5Qq/NGNoVgwZTXUitZTs+PoXGeeuQ
nLWubCyfs6HNBI0seLPwUEDFiEz6pQYwc/QwgNmObBmvh/5V6JEp9YqbGFRxoEMa
U4jvpjcKxO4v1XmQqRzz+VaHaxaYvdF7CfTnHJL4vCI3XkWdht7DcYhZPw5Gc/wz
twLX4VmrohynurUNOy9OqOoBDgpN2oYuEI2ldcqUzMn28r5Ntexk7ckOPDdEX3z3
Znv1q+7z8KEXSYsWlc/OmZeh288uSW5eu7qoUDGAV90wU+XrCtTZWIy6xxTr2L4m
2f7rnO9xj4fI0xec930m7w/bO/Vkf+n0fc3kzPzm4loF4C+rUV4aCezLVpK+AGy+
J+hf8E0neLNtXfXMuRlShYTtdFLBL39z/YNZhGvveSXuBoGflac/fdFlX3T9jg5Q
LtwvxmXFXDC4mmmCn5cljp1w6USJ3+VZ7bPEYKFWZidaazfg8wZppCtcZGsvPeB4
kjh3kE82FT5Ne47RNMn8fnzKukeN9jFTnrBjA3sAgk9fEVyN+mm5EJbdq9FnJMu5
Tb7qhfv5428ie+0ZX/+eFNr1zq8KxOjYRIwJU21wRh8Mw/hSJojN1qbXNWytDe80
DwUs2rSBpDh/4LCPQkut2HdQ2pH6x9Z8yeARP+GQgdqO0gJcq9cNZ2D/AqEJwZ/e
8qFsRJ9Ji7IPSTOyRs2r2bq3c0pQ8CvwH8EFAaCx05Relc8E4PO2EEbAWR9S7YZs
aPZ2yGj95kTJ4pw7etboMGbTgjt6cs+ShZ+uZ1dQbDYNQxbPQhUu5RJ2Hh5uMmYu
fieUlK7a1ATB0xAoT+ydj+XAUtAR/603yWTjGrVu32BVMokuqeRufbyXTpygI1DB
2P7u8ewj5xAAdwMmYnrI0AOW0gool61dP3mHOhg6fSQy+Z0oIXNSB5uNJcGES44+
TYDuV55e/wzBSV5U0hWFoIkj/a9TU9TQe/mpPB5uktQFbohYLsdSRJfiJX3zlNQz
2G3sFBOj3Ww4l7jCXeKaayE3T9APtDj6Vd6xkPSa9CLXEa3BlBD9LzDxwqkahHIS
tt7vSadS+kpQp/HNpxDtv0B+lVZ6NVSMwEXB1iC2HDDY1slDtJfLc/fDP5ooB2Ez
5AuOb1wq6wrFNPnWRH0UuHWfexE6OfddhLGhlVrEWqjTLUJSSyEYdCWhzQYl+jOD
q21ybJimzQ0UT9Ycj3id2ln2uGZNrq1NARdJ+ieH0jwFdvIMurXWyLQDl8CEnseD
0/jOYz2LtVcol7iegF70Eva2govzaT5PyMlgzA+lBGiRMoFqaGdc4RZuzt8M2yCR
zpedCJpq1G/FET5C0XHhLUHVy3Ue60ekw7bpqhh30F+MJgp3/cG3TYha8fPdBNrY
5ZCEy1AmBEsKO44eAJtGGu4u8esWve5UitF5y+Q3AF4dJlUOcJyoWfBLs62gqVbY
uLysaV/FDW6mdz/Ve/x0I3rqbVvRNV6RfZ2tgrxNgwPqq1NT0N0KU5JKR8ixffmb
c/9OAnaQ5Q3YV/J8wi4n3SsqEIexwDS5bDp5R82ZSOFUt/QokHi10KBxtg6KAKiD
HssCoVjOm2CRvpPMAQ/N3HsP+bweqtJSR0eJeVJjANWhqiDB9djBGVOYKICuVU3k
fRmFOIBBjMEZ6cIbV6itEZBBg17Wyq3wTFsO9OtG3VOkkY5i7MIcKqZwTPcyU9Bw
LqD32AbHZnQ+LXfmX6++WkErpBTTmnyyCkHngKkkseC9afx1vWnYNEJPLhpznXta
Igt8hfcG7UGBcXCniHqmd/ejUhpw0I4W2PlvMO+vKlFVMSNmb2pjVva3XSaeD6DW
tLQ+5pXMpiVdJNMSY4MF87avvNeu6Q+vNcj1ZhWsT4iV9zY+XYaqn2dqHk0JyLJf
jsQQ9lvHsZejt8uHS/beB9UVnP+PlzEUBTRKteE5UdnAw+/XytKWUiPpjwFQsAGM
KNwh9WslnicEWFsx/VKWES6GAsrLSNwx+j57cTmbkEqZzpdLaPyM1SsQDzjnoEGW
vta9MWqHB4fnSZikbqkYXBwQSy54bBwmV6wzyrRqhHjNuZlfL66690hxq6zvxkr+
b+Qkj3gJAm+AsWa5uSp15VP8i0kzA8jDc4Qog0hhNB7UZzP93YlyB1GvhWBpKHui
gqGdb+jjhHR2WZa3x7q2N0gXoxcs0pUfAmUTGXn1+gV2y2TTDVws4joFJVfEPVik
5kyv9d+3Ev26fl6n+dPR7M+bo+U+O8Tn6xVyWwzaiscrSv/RmGRwpFtGZtSCcWw5
ERrgD2FpufVGwzVxIaHUm4ypvTM24DRjjkq0BWD9qO4PHmi/Igj8sbR+g3PXvxU4
fmchBKPMsTvi+k3jq+dZ4HcO8FXNnZ7nt96PmQA5GGSsP02Cm/3R9k7NTuuRcx/m
I/KK7+ASJIreEOSQO9E5qFE11Hf2pCYR1uKb3yUzkYsbFnhqm6pmVCfnyYWVZOkT
a+849gIHj6PZYhq0a7ubOXUxOgq/99YQMb4ue9V4Cg5OFjNNQ0icio7w3bl0Xwym
Q4NVlvq8Iw/NXnfvC7UfjeF4CT1FhkoVLVA8w7ZS5pPKcS+tP8vsdw7+zCiazcMp
mSDUhcnrpvyuMwgmrBOZLL4l8yc+OE7wBhwCpkWwmsp0fvAML+NUEficiYBd2Fhl
yXWrZrrxcrC8ZOv6hO6SlpFWW5VzmSJcyjnmqXqNPFJf39y2A+uymmqR35HjJ5yb
c1cgNssNq+DsnF3IhkMZ142HZ+OjxZ5+MiESL3GOefZxxMytYlP2zQLzbmlPEOM4
YtWRGx4sgd4w4O4ldCKRiYZ3buZru0bcyyNWDvr2nilWLjGkHEFZtUPaTIjdaLPL
F7dDWwMDbeUQpK850eJeWVihdPfAqUunv2sY1v3wbOBjLXnlDqEuG6iMDxPIFQge
aDCZ4q2UfyqFn2FnnqfyM4kdzu3325Fe3/WXm0WEiey2/s6nB8xesNxd9bsDLUTa
PvkHiaMOEBo3r0/rSQFalH1iVjNfJfLbX6WYhpP07KvCmqITSPL8YqSD4o4Er9UK
PXodkLrcyUSlyXYyS4OuUZrRql4LBLLyeV916q5SboxlzS84zgtb9YR8Lk6xDpzT
IwcHVM00xV8E7DQ/3XRUixiyakAX5Omxv2EtSdrfCEO2EN1xsd0Nd33EvQ8PF/U6
ECdAiIDPan53i3ecUDBE+o8bwtNrmcuHPfvFgEZ8qjTFGSNqJVeatde49NpXuhZl
oK0y04PlfbDI+0MerZ75350MLkeAsQk5Ou8Z/3C9MOttOGOoseG8bPEWPpWTPTlB
BmZawGL8Fvx6deuwf/HRmMlLNTE0BnTSn/PU83v9QyHW158LShBipfv/Pr3LKRQ9
ao4I5+5U3JwIiLsFqXT2s10TJ3O0hWs1Tb/lm8BYDL0JDlH4zN0H+JrMRvjfYfLD
A6jph/cQa1n+J8CmQRPV5DYZ5BWbq/jrb6evZQxce3eGdKrq8oTbXnyPAA6KWuLE
G0z8BAAFVx8gUgjNiHnSjNCEHlk6CUnz69W9fvhGgb/VwlRwCG/aaJFSDF5BV2xs
JiSmhy9/Osn+xTRyvHPzHvDJ1/kQTyqh7Nrc6DPb+DfEt2gfuXQ6F2thkPvZTWpy
bbm0TrUOo2HlqJtKabcCIpq9eHhlOK9U3yTeR3gzJ7XRyowGTX6b7TKz054eYaKL
PNWYFTCesbhytZ8tsZvUmuwKW0waMSNQnCxR8F1ckWPWe4sWIYxPL8TvG+1uOW1J
7zsOAjzLr4daZXiltKHV6NcKXJaODN2joFD5etXW0Mn/9Rggua/qYWoXfOHIJMiJ
IkAJqwscvqjy+H4q2+ragMJSDfUGKKvdnp2LERPu/a2vR8iwqUJWtC1lyPT9tsgl
ziIVImPdQtjsx/WvBgwf7YF8ssddriWawk6eBqY7SerX+G03zCSDX8Enuc7b2/3t
KPHVmD7W4HA1DZbNyVffUkxJqbFLY/cDRUHGsFIhn6KDyyd5gIqxVCYyORe0Fuoo
+WUnUBsxBEbg7vpnkzNdoBEGoJu3Fr3M2Q14b7dbMLRgtPfwF9/s+aWDVmGq8Ilj
kLuR4GJB899QuBkbKn9P6K/MeVJdqvzS4SGaQ7gZCTXAtuVkCr0G11XGiZFXwMQN
VLIon9QnDQ8f/GjRYOvRSvMmzd5cdl+MH6v68x2nWVsOBJuR6hoGy5gM8/Ib6NY1
0a5j8Rc/Y/ZMrJxIH2Zu6r6bEysG/JRbnmRv1IaOrMK2CCqOPs9gNcOiSu3elICa
bl+5XgVjpV7cQSA5wFLHnnxi4jG2cd9+TZN7weSivPejMkA1dr9LvBCIfo6g6cWM
Sk1AuncSCXJpcDRKoH9xtFKEAdiBXJKQS1htREirZmCPo10GVG/++PPDA02hCxpq
hHKsg9lFPxZkaMsEr3EZzlJvapsYcgGnt9eBoWtMGaPH7Ddvpd9mSdrQ6SFjGuYJ
+0gMFcjZu+XJhnMKbXKaXHuvqw/30ujniVo810IWiN4K5DlI0BaFp4di5Iuf6Nz7
r/lHYPCi9F16vwatG4B3PA0/YqhTcQDA0qgabafmyd4vGHf180x1ky6PqG2kNiaN
a7fTv4F6l5ZL62VndesB+9CaFfmBq6hqB9hfgsuMCjRQjWmWxg+lmQtCjdCvAMA5
9C4gmqUQaz90C+OfLzzmlgh+xdcRiOEledyTzJwpXLAYUZ8OrqPx4S4X145tOJyQ
gZy0B6cDKYOJRt5G8QoRy/X5RiVMe/+H0o2Dw2Th608oTkmOMPMsPKzvHo36Yz4Y
KvKk1CsMigBQmH61NOETjtF2WFvPOV5YxWang5echZiDn3hRxxFLDjhCXF8mp6ED
7E+z6YcXfA3w9frAvniAro3+z4f/HS1V7rOuomJ+LN0DoozPXBUgpgJn/hF2DyHP
b61t0lf1GfYkvBA22yVNftKirLQ2LlYfr7X/TPw0urxwz0S6X54VqP9nSs8yy5XC
mv13ptN15EEXFmiNiwyPoCzg8quPrhM1hcfWkPvG+5pt2pXh2HPtXtoNnXG9QpnK
HHU/PY2H05WPjfYfCEywNh+wwQKeb/1Cx0qn8XsZ8nNtOKWhe3nA+ESTcXuJkmj0
csIVIGO0Hf8isQ9wkwK5Y5ZQ+ertEbaIJfoibJJ9PrSZa+sK1KvzClw6g0LMQscY
yFMdLyxYAu7fvKFT/UWHlwkAeedv2tpswfj7ulA0BpEiBn/qMNJlbs4BFvrszxH4
4f/VRCKI8KR73SU5siHn/zoXo53JsRQJSwRCcXNqLWLa9F0xx+pDlfxqwO/B3bfx
XPiTstKuyzxMROCNpqwSs9lJ6Ahjpkqa/CPlpgwGFgatVnkuJLMo71+bTzQybHrv
LyTaWy/IExHZR6sOqzuHZ7gTt+BclnZ4DejvEPWAs8xjylqMg9lhySlRiK6UlBUm
uFBrCPiWdGPc+tkIhWBFwZgRadVVclasRXSah4BY/0cT1hjhm1SR+kP/417flPFX
8REpsxTAbUQ50hwef2XlbfJj/7jF8J5hnzgybmSwWyXIjP1EBT2+15mJEGAZO5gy
hhAszUiI9hlPdxnqainfRR/WTHVVauSavHDQ6FOFENVAikDM3BUduFkkkxsw/T/t
1mMAyi8NJfvZdbOUWPKPC7/K9ROw9GLNy1PGyF2JHkQNckFltJRTaxQeaHyqpQC9
gMMyUkJpNMYqSZfbOi8mZJgeju5SlqNN1JQvttLWJkchA8rTXIX8TrkR8Qt6IXoB
lzyKkYSb8lQWc3uFIGYL5rqKtMTOdfjwU/q06gj7tIrO9P3YO5/usZ0aElhrpf4O
I1pgQSLamtXe4lTkKRe9wIMwFNMZZ8kmrtbvTKMVgnkzjb7XAeNDl1Oy4T/fA/+G
dLwlQRY/AveQw826yfTxVAShEFJI8YkHMmbuj3dps0FF2INIeUwYCkf6ZN4hvA8Q
MzfzkF66S2PFkM++ood9o62N88QWvnj1MbDupX8sqlVz1aelduRd700kEf1V5ww2
EOD30p9DQg/q8s/OYXWgVtuzic1JMZcoWyTXG1oYe1wfyoZhRl1fYnhIawpdxmFy
jnqcQd0Z9u6vUpKucU/OYRVb4EwS6vc5SwksCveKAtluRGBcFWK1HYJS8y+PSBqI
DDEIHtdvedgfzb0lOmyN9mpxVne4Kor2IHdEuQGx7Qll87VTRPVqGAMapzZ9B6Ma
w9tDKgTg5p66g2XUWyTn24pcHUQNwIc9Zw0HbR4f0Q6Zu0IPEvDC//iBcEoviUTJ
JQq3dr35jRjxlGdQu16mrFo6A7cOyBQm6x+SWanX5+IXvTc81yk1pZsd82XpCg3N
FkNoKN45EJBWey47GURrdfmHH4rhPMXboBDuP4iDCrTElfZ/w6Cd/NI26fhfciCo
G2f3BsKmzIH/3MatZ0fu6cRWWiRTTDZzBhqLeCdhZgvuBBDhE+RVw4f0IvoRXNJl
5yd8IW0jQoFXAmdARBFHAHO7nl/eFHi4b2+TErRsZXi4zhBOskJZVwf21mKqXCdi
yYosC9moaeFcXwC6TfUYKKLFB5QWN04Nk1D4pcLhwYRUhYvOX5ywGF+4PFlUdE1r
2MsZpuDupqrCnqSXtU+dIAa7oSAsQxOpk0MR8dPrvUiL7wnFsyFUkHU+xL7Qvxaj
dFayqC3mn3fGy5ojjatu7grQQjA23zPhfhUCLNdc6ZAb7COQtdUq6EbNuvDMmuM7
szuPN70mDbfwDeJ/O6EMbl0ysDqW8FdXtT06rHcKNRsoWGvZrLbKMGoN6m5e4j+T
jaILk0T8bFKZtaBObUiqVsoSzUwWAezGixnfJh0NUaQvNxZJ6LmUXHrg4ncBlOoh
g9XumK8Qb1iIo9gVG8ZP00nOnlcWwVURhhqoQ1SKn+7k4jnvs3ACGlaacwo7bOTT
yCH/lZrJJ7pleRNKJv1UKG5cGJhnsttOj6G/Mu8sGZ/4dkQKbEOJT6ITlHIZnTO2
uRpvbZideaw+KWPt3DrHXk//MYxaYTOOKV0Q60CQYjiLcaKlD0S9JHHf7IkFaVfM
G2VE5HLt8t/80IkjYGuYu/BaaLNqDbvc7r5DKjV/4GCprOGP18/YNYrl0iJJdBZf
+/4btsS/he3CWe1WRCgEBoMwdJV/Bw+NSdr07VWbl/GdyElSx8DMeji/YpfYc1mb
TkUn0UOK+tKBsJjYIvQzSHSFh1vojDSbmktk0IrGie0vx93jz6xE1Bt52KEjzRAz
FtfyxvsE4OZ/sUQJ7j71SJRb6jhA1DnVMETWF/e2Dntg34MjiesIHL/c9NXohDMW
1ldlOOFdpsirC8gEygfkAwHI31PpZMf1Q/WYPgzNEjfr6FSsOjJPz7MMt/sHLdaQ
NgJsWGKQ2W7BUZ87RwULZft/aSlqX8vt04Yu4BaCD0sSfijYlmHHEBEZ26iAUCWj
ggko0eQnoqOG8b6ig38YG2ewNqy7Oj1dY+5cCZ9vuVMjmCCdN1fUfEXe9fyQ3PE/
IzvDElyxb3alolmWckq9hESaO7IgokEefdya/RXA+KPCe+p1jhyTAGc8uJsDOV7E
MJI3T46EvoiEXETKS7p9+0iPTqViJx4R34UTiSEzJIOQpSRl0aKDYnOzqvpKeOKy
I+itD7+s+CA7yyXz90aXl7Asw4kKPlRvAaR3yH8wciJUB14vcpj4s45XqrMel1AT
3fArDrdWV/ItLidgGKpyAuPDp0TG44Z1rMNmmG88/VUIEMUiulZgQ8r1wbr4aFEq
kfYkNbqkFy2nVgM/hE9Jwq50HkIBbpTMahtMwGydY3oF6suckjPt3xvsGs+Cf8x8
mFrS73F/zjUNjU/UIY4mO3WyJONDCYVkElEpsle11q+btnenZVuVsSMVzLgpf4Zr
ZmR9/TJNDKI3aQe4AU0aD6z17LzHyrkYf/JrDi6ZGrwoG+XKmeBwxWjRuyTBH5bK
wlM7RVdW/v+u5Tsj43I+jY6AhsQKyN2un+tyC4oV868Pzwh0fr4RvUnRUK8opk+C
c2kz2brcW6A8T3jqTePpcZgggW+2YUiqu6acczo92nNwrNVgVCSB6+iss4BkopiV
MyxWGkSh/hBiXvytK0s4YC8deeJ/YgZKKLzF0C4jGcc18B9MT3KVfTfuidfy/q+R
bwXVw7pGyeU1OceQhqZGYDpdxSkDc/cMQxq3Q70Dna7N9rW10acx4dHd9BdLgRFt
k9O4C7B3psIf6RaQxR9QLAGu4/cT5HqFoi9zqInkuc2WsNR9Qv/VCRLx0XlMII9T
XO2swVGdBsLzfwjLlCUFAw+t7HdOJLxyiLmKeTMGlV0tz+Z3DsPWXHudGascZIlu
QFqLs2Od8Ji7JWCxSuZQ6bH/Two4/60hQFFRc4bcEMaMBpgQsj4jX92yiRF4Qjhp
2l2/kTIuQUq0NNdoCumupprn2LPmmr6APxx+wB9sxJhWQk7mY5VmdnGqfGuMRaRy
zsVvnI6PImnzWVtJoRqkZOIM6NVnfyNk9CZKZPcVPntrH8RoiDnk9TXtjcZqR/Xy
82nKKSLJXzAPoQF1sdULRbECcOb31rGCWkEn+ZHsqKI3N0YwonaanIfGlxVdBQJb
C8zXtNF6N1nMGc3ioQEj8nsKUon+kIVRMKSFAuIeEpcJ1cCbYGvG4A0ZKirOvA9s
gOXHZ+8oBlbIneXh+cL0FNTfo5jHmeJcSedm9EYe+z8Yfwz/E/WzGc9OpimCSu72
VowlC8i4QeGHs4r4h0ps82SS/egbHXqeXgF6O6+7zzJw3B+i445z/jPDszNFuNCn
9R8O1/v306S6nxS3K+BTR/fo035tFbuKzms664Zxt1esgAib47iurYKA7LOwSvrQ
F+GgGl/y0I5YpxWKYO7xmCiWgP6ZbPx1kBZULdFlLmwAsrLsfvqDDLtxCofJ+IHQ
SvSw0t7xemv2i/NJ6qult7fgo2HU1+OslIeF0ER+oxlz2BDTJ1J3FMlCgYCL92tc
pRNGlpWKgNtF2zzX3F4X6f/JfH1sGDBeiCNiJOpLgtkssq9FPawMaP5vWLtIdQa2
aCtkv+yZitlt0LrkFToe/BJW7ZAK3yXer+M17quxhysVBcy3io97fpKQdbMD2o4O
+NN5b22x+SUnwJT+gZ9ynA+q56aQTk0fQVoVzgduraghRKvcCl9Z4K1IRx6WNrO8
5pAqTNjS0K6mVO9E10WiBksaSBYMwLWCq64uonb8851V8t618Kn64rPk8/ucvjwm
NDtHrJCBMbZDD6ls9gPT7pUAQrz7tv9y+a74D7RbfGrOsUemmdWQRyaczspHwefQ
MJnEKJapuBSD1vUkNVsqkhSR8RbLvjPqFCs7wafIZ4dkuADldm1THuYzViyBM5Hm
lDk2wlKYlxCE8jTHSHPsXYczRKVrc05WL954is5SWpFIhwyv1aZsN7vKklNeZQTM
RYhgOwQQP4dTxJAsRa1lppPV14uB5PRjSxzw4vl4U8uChLZjScY03KdYuSKBCceN
fMmeePyLfFPFetNTTov3rI3ILFjJgJC6uMdu/7cDa8VE6RKQrLl7WqpXKPULYWkA
HZyjHfX2llRbZ8GFGGMXAg6Qid0GYmEHcCiPAm0NLWKzCt2NsFb7Ez+3fgKWHefN
P2crB6c4ly5IZ5CSMzpGie+GA4QdVnYotyaNAYx5UylkYG1DSMM0G5D+PdPQ4hHl
e+Zc8xIV3S8UDEwmMy8T2QXX/lqu8R6Mw8UKIraJbPZtGFYLacX1ZlwsCM5cTlQG
+ED2nNKD24aXcmdAk3zgA/RmyXdVWaFFezNynrWgDGBmnDaQ1zPxc2K+Z0qIKSQb
E+L9ntMwjb45QqSvK0k/6OZVtNctWRVUURQaQawuVoMCwT8e8z6E//SE00v1P+jB
JiOCE6TtPi7Xc+VnpeVxbHI/T0JW/kgjQowbpN693XRQqit5uB7BjnstqBxUzuku
/gSXRfXpQ4FN4NTc5rJY1W5h++UXx7yobNQ7JtOwxmqf2xgicJF/e3UuX020YBd7
okrodFytdkiIdcdQUVRDhJP68XDQXa6IGrNxhL105qgVXTHTQpN0i49758n1adnG
wZz9Sdyo1pctJjsyIV+3ZUHQIDcgF7znykKMPBhTTubpAyohgMvIFHGst1mTsiUc
zAMvF3ioAWOtfXee6dzyiKi6AnDiLdoe0rxL6FowTI2H3pxyOYLshQNchqeHLAZX
3gqP08fgIj7Y6HGJ+XQ9zU8UkO+uGWOetqxOX+e2Z3CM1YT0HX4s0yv/P0omlDZ1
I3Tbv6YzOAK29qU63dp9FEXNTtoyI47lJZ7nTHwvk9Gpu8MYiiQ/odFjIMVW9VUm
AJxormuRx27qOojI01MMD20naW1Xm6XwFCrtuuJXXeu/rlGnkA3DFxZeLFbfSEvf
gSJWRxd0crE7PuKgA1LUOpsHD1ht8I65kToDS7TcNjyeNQtOjemrocaQMgpmtr4c
k3ChZW1RY2DVci2VUmC3er96Uzrsf47RJZ+RiVUSIYEC5aLHvq3sFL5ARSvK5kdf
aZwbkzoRSgnV7MsGGZtaWIklVEv9JMrgVGrPIWK3DwHCqTzikS4vzZhXoW5SWXby
64cfb41urKmIBoueneaS7hWsOl5+JfmBibJo5Po3wS68OiAtxKgn0cyozsf+P0J3
q23R2rHphaIcYW4hS8gg9pIgwGup76+aCHPcVhtygiNhUJscBKi9kVHfNmkKph72
bww02ohxjBaUJOMvffzxvsNNY0jqLA84v7rKjafa4xk2qg0SiBqQ1KvCfiyjyVPm
ky5G7MwZlXHNMP7L5P4KwyQaPWQFAowTbYsvRhyhesDfh9OZFnD3Zqt/T3g4WlK6
jF0JhrmKIQ4soYxneYfcqVv7NJbXapvzHF4TPiM0xoP4XRabB9yaQrupyuT6Xy4C
3tKxJcXrcNIdXnYpuQPjvuTiU6aj9GJsDxZVjZuAvWpK8Yj2kvYp8Iew7685cZMw
3jyUe5763t+l10AZ1TbmCVVJWgFXJF7eVlrKJBLnu/WfPx/WPerNhVbiuJtbgI2Q
IRsxTmZc8IT3yloeafOlSgZT+8xYMaNDXJ9qbRhyfD7ej5Ld8T2oyRTiGIn3dqpN
Cv/LTjTOp45zD5hdZYJXH7mwEdjXOZ3XIJNTEWEHU02K27IN52PA5x1h1q1mnQG+
beAwJ/KNIOEwVUI6+I4LzKrj5nCNfi8mgp6P83QobD6rt060Ckgv5hFHJANt6J6D
6FPkiqLGpedqL0QlF1lgcKTy/54JIs/Mhr/G2dAQ56S6K5ES2FS1QRIRnsV61PJV
R+XVPTGQP1CFMoJDtfeF7gcY3NYF5qDZDyyzoSRdWvMFdsNmb3firlnJmI+9c3oy
wrzKU6YnZaj/nFmkpY4xpA0g2QRG2qidHClvxsFeqgcbXf4LQA7bznkt3bvSCV/X
8ZjKml99zR0ZkBi2a9BZF8VMCFKM2GYpJsJqeUdsqgnC3DiCqmNDmzib4DxWxQZZ
wF50kY2PGOfyIXIFaiZMBEU/YefggeTQAJ0Lhnj5I4FD2mA/MH8HoVMnLjcNaFiy
FIyEa5+qCXJ+cJHt4+Y/S8BUpgS/KjlQHSL8wes089xZdahaK+QXc9ph5h+Lvrtr
NMl9YKOPdOvkVo3KkYs5QFDysSt6RzLFU6dMUIOrr7HUcIIPEsI3AejYp8qN6BiB
1Klv1F0sgScqzZa7gVSzij0Nf5KDw9dFHpaC4Xfuy7xBgwVdklblkjvf4fy2XTtU
46vTXwGLyQavMia9D70mJYL/npjl4NqGuXPm5pj1TFmlVXvgZau6NabPrBZR3iwO
ZXqoUvJY8hx/Nhp61k5DiAc5saf5xqvE3o1VFWOejreAe6EX7gajc9/SoCnIvnbn
tI9aLgNQzSYyzBvB6FrVp2Eq1My/kb19zZChnTwp7l1VOaF592ma98KZuTYR3zvS
x8HCq2jOOXYAIwuf+w1p96VK4jQxGBidV+QvwqsvO3LURsk3ywgN9jbm1fNZgPOp
rYJH65DCs+UpctKGkA1TyahBJeIDhzTlAhkWCcyvF7KQfJLUaHttbR8oWFUChSVs
d4DLthcTycxR9A8ZNH448GW7oTzSUJkyjicjanxYAddkeIo1XD7LIuYOyIB5/5KQ
ls8l6lw0wZwfofJ8aoncSo3XXrIKTpno5uAVx0Tpq1WoBm/9B7w7DCkQgR8u2VJu
52vABelXOoyiGpIbA98OtOUe4mzEkFor18urMxTHHTugKC8NaUFY+QyKrJfMU7m6
I/g1Sh4yX58eeDsPFgGCOy0LqPdFE1dC+7qjOFfOhvelxQH2glMI1wpN3zGbOoPa
o6CHTBGhg3FwHqBsdx65rweqPoNGPalq3Cz4E2J3moQ/Z5qAcYlpZ1qhhfdJA+Ak
m+4M5bHkhwRW0EnitXPB+15DF4blU/73uXjXIguwmqgJ8DDiHMN24C+0X6iM4A60
YjkrvQ/9k6q82pSHbCa/JQuSMWgbr1WiAcUUjUXqsuSoL7zBMGYG0F7o1GP87OmT
C8aLcov7RefBK9+Qkp2IICLa/bAJqkUdfCy+BU2s2LqU+b0zsjPt9P1xcxzvzWM2
1N043X/KEdpUzjIc9iEUzAG3CZxfaqOV4bSYdVyBFwyMaWUnNjLAO5N6smZufBRG
HFbRU0AxmknQ634dOmZLSIjMbpg+SNMgGlJzrBFMBFriz6+L4Torhd+f1tAxg+rG
HzDvCt3Z+GbHcHlWGpLIkgDbslkTUQnZIGWP6dpBOMdvG3lg/olkIEtWE0e3xocR
qmCsg0GIeEnKQboOdV6iQYRxgNDoCMj5TlBr0+Wq8kMbeUOwiA2qx9rSRUmqylSC
83mZRuTYGfUZvKeT/2SYL/Bk/O6xtpJc+f5vndR4cAjiTXGmDGbIpjbN9PD3kH2O
Rwho66hDN2eTMbUueHqDM5KIVmXsHeeEwb6c7FXMkOAj9HbLUHM9Cv68Oim163ow
ZEYGMr+9ZxhUIUfAz5648D2aceHAjeZaHcns8mwdEsVncMl55j1LejTN9y8Sm5Vb
ox/CqKY4oMSiTpFV/onwG6jjFxq7korHdLpgcmYa0+b0Z/+f1vYpauV7XV0BcZh6
cxaZdE+l10BzUxpyWibIjGFVpD/SetBg4EMvlljCl9a0eALrWjXfnRkVPwwTQlOZ
APUAM9I1O+7rOeE21JOlNyuPP9Ho9ZG0Mkgz7q7dQ4LPd4MmkR3QuftlAlWzE01v
cdHDmPxvsNq5tE2Z8cG+K1nVbzsDhJAtRekelAkt7PhHHmG/jlJcTOIGcktHn0Rb
QMhhWAjIi6Ta6bo6nsl4kJZ1uyTFaQRcmg2Ai4pTgFGuq0vAQjxCY0NAFVKN1c58
OJNOK+EHF6GHz6hfKKcSRoYtbI+E99SI6pYeb6OE3y6wbg8WBSwis3Y9vlhUVDYS
kGuQmF3H3d8/5xDLQCsWXY9ySWX/Y7gz0nl5iMO93if/WAV+BMhwjMNuRUX9Abm4
8BKii4+fpcM3N7oQl5k9S+cDfdRBmDTvwHayYYMI80K7KQalXlEu36ijmmH9yXyx
PculY3uVOHLS3b45D1IhYmOj+PvS29pCCCxfjpc64PLWxXYGQBLcmAIqFhgbkQkc
CSMUzUzhxpWDDsWb6vyb9D1eCsAuye/h3rADj1mrMXLJS5bu4hgcOrIWSvGI9VFx
PFf+Hrh76ADpU15/UvMWsBNzhE1ZX9aG3lHoiUcW95Yu+HQnthLjGz2bbdAwOGDw
nNFpV6DwORN4481HKUMxQ3bd8Gs3s3IvD3UUTdT3HnnnLiSvzGMlp7E9U2hA7kwI
9DQehfFOcTwhCuinRzgXEaXwF6DNoHIxHJBbDkCbN1xcEEH/+J+otQ5gXaHO7YDg
M+cFvRm9ezI9AQ1mrzUKyRwYglYIzRIHq68OXdtCv+/InqdCugZLM5FcpHcegWNt
zLdCnhOFKePxN+44WSua2XKy2ld1Af0JlfRcT9EwKqLju2CCgLOTwbCzzjLzp5rA
kT6F3q5ZLqOg0uWDdEw3Kp0nGfS5fgiscDs05uGjblWL9h2LWxE5iJVPqgkIQI26
clWcekjHGHu923RaHNo2IeXP/DyHtsyunevOAAjt93LyoAvE7ofBWbtgoN6ax7Rm
sKdIp5heHJi9/CNnCVrQC32EsNGZt9H+DH8ZgH+15rh8a14IC9fdcCHi1cObzTDW
bKHCk5jlOuZ36Z0MljFsL1N/HbMxagkam3CxTaKkeDSE0Xg98FScH+DXdoW/32rP
pi6Eu2oB4YGC26T37HSPMUqQwwLGwVzvUjJCFq7P+aBa0TMhgYa98/enaWUN1Gsz
I+FL1XXBrhK3kXCf3silGaHzXd9R7lHqKNwtoHuCq+DjdQz+wHeY2UXZ1DXhFlJi
sRVi0u10M+SOk5YpuNRBGEXOXkXyvtyjNjZDhr/n/+m6A+M2razegqWyxclWvJmJ
/VnFecWemiRWkhAqXJ8RDcOV7hGDQpVb302kHwlcX2c9MXvdrPeeH6cVgai5Oik5
pLadFkxGSye6QfrIGcTLfeNaPP+FADXCHyQck68hJScsWz79BlYKQyox1FxWqQsl
W3qsks2m5W4mVwvsJDRLYOL/CwA6ofFzbiTY1bhcpiorbOUsi3sQg4LuZ7aOMB3g
DCMwNlpvBTn1mBcg6B0S62Q5kceVD7qKoy4RiZwqBfJx70hkm6KHFOyfCgDXgCiE
XwD/P1pJ4OBTIY/bp792J9JNTRwyXwnpIuA/JcqBSQgBXQjnBHskrxl/KwQUwGM+
rZiEfkLI5NqUrF9YqLyB9xmM68TwkSGFfA/1OHb1K8Z+hrcI2pdfOXe8iv/tyf/n
UdviXsG5RfRUjqWfayZxftShltci1Xb61ebNLjDc095lpDmpwtd3b3XJ9nzMzr8m
Gm4H7RFI6SqkseKT/KV9yLn7wpA96fZXut8z6N6hYmrVy6Sm1CG7VLpmawmGUKzx
AO70yWLu5pJfa0QkpJxlWbg2eqmxYDLTD90qIpZ/B7hbdBSqK5oIhK1etgwkMgcv
IdzTQh6uVn+2/9joEuSJDoSu+BBk40MK9foHOr8Dft9BhTPpzD7wGnv1QrJ7HLD+
vnTBBn7jeqQp9KfXyWl/YKLrILThCLQYzvb0BEWy6FQ1lrnnL8mbccew6LFsth0+
eJer3X6vmWO/qrdDyOkOTZg12mMfTGMlJFvvZiYfsu0JLuGa8Mwb1f2gU4WIbsni
4H9yeovg5juLN6PQckK+N+Dv253f7aa/3NXg9ff+2xL4ab4LiYJyr82yXGBhw93z
MmFGk1+FIcncR5WfOLeHy6cSdbM1/qJUfAHGL70zDtjaGIE/iVs7wTzaQrsoflMq
GI4VJXos3XjLY3Xp44dLKOG1lqRjuNPOpjqx2+iUUyIOLkrMuyPV7Hp7XjxB7ep2
b6E7ni7BC2MJzogalerskBo+vX5ts45KzBDgYgQWEhBfzNeJfF34qv3VbJdIzter
SB/ceZ0eIauhHgNlf9sO2mXjCtFc+BPO7UCVHtb7GSRt6caXrWglmxUXN1+ntiaO
MxdHjXINYz8rdgs+zkGeUThwv6vNOylZcZDztjbE7I2Zc1u5bKqfcu5+cRVGg8Pj
M4BcwtGkj/EeJ1DrvDk/4ruFz3/kbl19qkaCWEcB9MyVpWBRdPfQtPjXospdrtT2
9sAH8GBDhvOj8ZDvokCLI7nwaAB6LXDq8xOsIx4JG5eEAznz+UXMJrNPqeXHqJr4
CAqq2FBhSGaRQvdspxW2WqnZsqGR+hkd29Lqy5UkNHxvK+T5gWOeqVtKAQMeNnOp
5FtT/utPoBgnCCJy1asP4af9LiWXo7nXYLN/lamcZqGhiVCttSdD20ZtHf/0P/f+
bmdVge1F72hEJvj49a3rSsDCxoKFtjBicH8TA0nosBcn5/jDlEE/0lmgbUHVeamM
V881gZY14KNkyYrG+cyudkHJtwS1L69UUI2+9C5l46J6z+KHe3pozH7mCK8tfHFK
Yhg+1+4aD7zOBSY/Llu4g7Co1nfMCBUUGALgDLvi1Y0TzohvkckaTcfUi8Bc4Amf
FFLmeEjX4PCxGeTvdfo7Oznlrd6IzhkdCqK+wstD59gwuQeqQGBKzNWGaFh6HcUf
80FxwL+tEY0J7NvZZxD51xM/JKwPKJowXBP6+hU7avDMINlLYgDJ2dIgYZh5j9r0
HhegSc+NBGrdhudrl0n/2kqB9N75yF5oJtUQKd74whjT4ZUcrkQJD1t7NZH9St4M
WDYh9RjmdkuA6HDPhbu/WhqBp5mnaDeoBCr7jxsJs2eOMsflAaGWHPvCeQLlyVXg
HdK4XXzdF8xyQy3MmVaegVihDZeQjrbS/uHNE1iRUU5oW6Et4h+gLIHQrANMb2X6
Tkl6zzMcPJ2XjiVoQMjCssyLsUhpYVssfmeTg0IBjLUGluPGJDZ3C209D2egha95
SUzbdPxDdlhfLAheBRz31AIh7DZBSH2xJQ31L9nN5NpwyHN30J+TyRj8kwxV2V6X
4Rh+WJHyoJoRfrNzjx2aMtaJmBdb8nad9/KaircvfmVjMiLAV33KLFLbj9KhAWyj
35EBlswiShtGlAqHN0fk/IYv+p/QYISt18ojs6fu7cqgozhkcsoPVC7gbEco+Oy7
adT/Mat/8LpYaJu9i5BW/V8DOpSA6YzXHoVeOfhsYFMksjSB11/Z9Ytk97b8O39y
+HGGET0qziG6qTsLlX7YT6lX8wbMnCEcvrzGFM1SravpcUXXWfGtR4MmR8VVHCcn
7HEtShOeWKFE/G/U4eoTot2Nt6V+57/1uF/SeKgIo3Ck2StHccbfJCubY3plfs9f
KwpqCfO/CUYVhUzgMApGJuKou8AsnLUbrMSZdD/kiB2EqEkfuaADXw1OlYQ8bLfv
urCVIZ8UbbW4TzZq1zrrCuye0aaSi3Fmdd1d+65M/111LOf/9DYgj845Ut9StoUk
yIuGIO5cv7Dp9nW1WDC8u4uQMmpIbkqcfA8+Rew/X7zXwKmIkXpmn2ljdyqIHDlC
rQHoB2seL/+nip+kxU/IlHvTPkpIgY5f1QL/Yy3IGjGkhuRNSMTY8SACxVE1AM0H
SJyRN4269DcAD/AosT3cfr0lxvnpipIUbo0OkuVQfd7zWg3j8jt0tN26/+NMXEhe
Fu5aYUiO9Gpzg8HQbkIWYBsnW9VUsdISKyBGyplL5bAPOgv5YLHq/EL3IrRWGiWx
TQzd83s2bvX2lkLQFYGl+gqpnxRA22ouOkDIPvtJGYNwBQytD2d0MVFoStTAJ6Zw
G2xO3nXoqvyze7GXgZqNuz/aTwipKryNBt7fNfEboTKATbgDTPe+4PGRPa+uQhB2
EYWytTqt3LGdKhvWakwnzBPRZ0DYwqiE1STATmqIB+pfRdv95erYkgiBmdIz7xQk
3if+9TMAmcSpD+Tlw80dMkGeaYSWAN0AXfoW/zArY2vlCjfAUnppCMwE00erHYPi
WA/YaEHKgPkEw/MV/0YAO9wItCj/My1HtlEY1oplpt56DN8v8jK0qwAzCEuQgBLP
XnLbLS3NOOUl5peKNH06IoIBhi+QjfpZNZ6uYq8OA5xBpRiAXt27odid1Vb1/TGN
zJLC5oprf4/qFa4Qj2M+qkrUUnXGqhAdSefGXSSco5CwmkCk/ZHvzrTZQ39wCTpa
U3v/JsHuSpEXnQkLL4OHJYGZ3Ziv8+K2bIJ1MwwY+SQ20nKtfDPV9oXiL6zAR5vB
FNAbAzVjOehvfYoxNuBi2SdVVv9gML24qBcYQryQ10qUevLADTTQe2zVdC16MN2H
ecUluOwZg5x6fB3sWqCA1Z+wCPsb4QiFaIc3qf0MvOB+QJ6PautsJia9yT0PcDHk
o4bP/UWma2OoZ96KpPS3FI+gYs8PA653ZlBelfePrAHoyGsJ43uN4PY7gB/B8+5G
9bFCUOwddnK/8kAlixnHa1h7hLTf02Y6ElE22NDNHTsVkl5bJIHv4RyqevXK9aZm
iqcDXdnplDZ00zMj5QMA78d56LzM/hv/ek1t4FbdyanlhX6urTHWkYWsbLbRl4Km
GCLoTvBRjodwuoT/pKw8rv2Y0ISyJaKPwnGg7Aj3S9PTWq6tDSFAX6QJOiIftDw2
odEO0kl4h1lufH/KWRIm4BOvxIMLMZ/kXJdT6i/FRKCsH6kspDofExnJXoEOxuuz
1p0p9nmTd3osMsLIeDJE8zMF2y6V4K0a9/InOc3HX/H37O2O2mrSiLMMeE43G4HI
ssuUUN2ka1xqny45RR9ytOixkLWzLDglsLicrlM14hwDI0ymETAKg6u8X0ozdCkM
6r0N0T2jJdKnKNDbidHrQzGZmeP+AYMKTIvhz3t5kie9PVi+CX/a3XIXJ4lhBQyT
3akLfDfC0CqZi4fJwkr/tJ04aUf/ma/gJQIUrPLBLSaonvlBs7NhLvlYDrDFa1Dt
FV4p0Bfiq1gbKdIOQAngJgGfLc+5FE10N+2N5TZW0lOiSeUgViJqUMxhOKxyo6C6
04LQ3tEwnRjXK5aQzb6Td/ywABfwo24RxnvO36MRyaeX1kXXjofpnyaKYtstoBCL
Ccz2A8a9BGC0kbruEU/7xliq5AeF+g8rBQHKeZvC3ILlJsppLh3vojVXA5zpgT6A
5HJ0IEJPDfV96ld/7/8hR8kpICGR9HTO6H4JW+OKnJpFIgpHi/sq6D14LWpp8UL+
hGXZ2T1//LcbGkfIXOo7Z3CYWEyKQ6tKWD3Lmg1EH6Tw7wstNWo4kYSUSWABGpoW
sop2MudDTLfdicYeIZprsM4EiG9OsBHr9GLWnpU0kJr1BYuUhmuV9+bM/ev0suCm
UCBp/KjRZk2l+fSh6x+LijswLmM+X4V2OufvJ3+lJ1Q4T3rY97fZ1q1ezy9D4CrI
As5kGl6cbAeftb/uaCKCHv8slPyWJWlMC6vAzHVqWav/91MmHN271+b1k/Cz9CG/
s3IEXH4p/FEaqofkYEIm8lhi7u14p6ZObfS8zmRHmEkyDUP5GIqF/oSlKLsCA4nC
yk9jQ2ei6onRWHKhkPLQaKqt5ijtl69v8tfz3/jUzI+pkh2bbOLm0Qq0Ft0VTKHD
Zr7po7aSNCIfv9nS3X4hdFEqKS0YnPZNEHcAtHnaZVqiqoiQU3QEsf+7ZOMd4iMG
kbjXaziVUETl8pI2N2atrupHo0y99kULyweGzNkzsR56XN8VSiunnCZZS9T9qOMm
x0K8eB33Cj3R0i88PsEL+GAZYZnlTllLv1gDLscwkS7tnWsISFkzu0GcVsP92OHD
bElzc3HLoWEvmdkphLnEuBLjrkdJSR0V558L7ftMmxx3R7q/F9xCjGttWzCGPQKh
RdA7qHZLpTv5Alun5+WOZlUAl+vkqdrhsRJ3DwU5+7CFZttoLCHSqpByY7Ca80eF
n3KQSfYZrwU3qH81VFLRKSOi4nGTXFHxk4xWKMfYpoFpSyACyf99g6VUamADNgw+
9ExI+uS1jgH/0MjkoesA8N04PIyehHhdLgBKtYWvPnAfZa/ocnKSS1Benj/J649u
zc7ubdo6y1YduLpWJtRjeAV6J1io8bHY1Afy6bGwjbkiqqGXg/w+A/2MZz6bA2uH
e3s8hhryOB2SiKWsdKVyGutWGM5OJMMN4NjKF1z/Aqkbw3y1AZfnKFfxBpBav+Nm
aCiRYIUXb0iRJ6bqn0bsXfCYgaMhAKOTWW7gcC/Xp7yfGVs3oUfX9iAitGIN3wxn
ijn/1QWtDqlXu8CPTeTolBlaIQXWcJs/SQzuyd+HHwzEysA/3J/D/L+63BWGonk4
F2V3vJJc8nofm7yuKkGcVheQNoawTrZrQCZHp2dSzdwYMjAKwXipTue3sQ2Uy6A7
d/Ur5YURgUUYQY3hJQsFF5Utom0xB/JTWy9p/O4D53cnZMGCqO2UWFEprqsPnyTF
EXgnRcDSf8THubZuI5JU33N6OZ94ttg8OvbaQxfPX4prR/JeOCx8oZhzrJ10bFB+
XxOi6q6bO4iikHdLJAIcUA8yFn/F7aiJ8m0vrTefr6NNBIZe7ZfcgqLsXSfZ3Qj+
R+lqz5Bll4dta2kNf73oshW821dmaRSMCy7hfue4s+y2MHVgFBWBAEDRtQqjcknB
JHqdF/Ou306lc6yLBNMke8zGT65X8j99PhNkZ9OA0bhc2gbT9h+dfoQET3tn5WHK
dghVdl6M2jEXySnHMHt0Jau0CxNCBZO6m12V34zcevfke96WNzr0DxR67yBeon9a
Ou1W6Fv8m44XtiFBise6C6feai9OOsWgWr8d32oU0EKATJU5349DvtkiRVsJClkk
ewMR0Gen8nifJy13hRcGXFhIkG/YPNniPA3sA+NAoBoxI0LVimrivYOny5qrwB8Z
DVp38h6rWjHbr6nPMoSm7qm83oaDsoMSDSOpOIdMbMnxn9MZ+Si2V+B3ZXASp69n
ilayR81lRJYh3N5nHGWgn4bZs9OkOqBKfugykeKJyIP8ydnt8XQ5NR9HqxE2JK+5
RzpIDhtoGpRrotGmjY971H+K4WRdLUCtTmOaL0fQKvtNe7UTB+oYZxlhdU49R8mC
X1IIdZClGhRi65VPXVXFOHt2EAraRWfw3zF+RDB2LaAShOLdBJ/PtaM7xkY2r8zp
ERITCB7mjg4FksFBFG8bi/vKfUG/G/v78+YMjuwZGmkMgBPmkyC8K74BJG9qmrqQ
di1mxzLHZgItwk5fD6Hp/UF6g/6ds0RUgxSLtuZDii9X21JmeuTqYxK0upn0Twax
W9ZIXp66wguvfME/Fj+vj9bm4Ix8v5ndvP0hAxLZ6NNYDffgIwJPApYh4hiAiZZh
xfi6h8nhG8GqcTSBP0podC2rQf90oJPG0z5Z2XM+QtjxZkccXHBZco0K3eaMo5rq
oCFAOhsKrWGsR21Wi4uMpatJIKy+OHH7F7PcVDlgmZqQH9MLsyEqh7QA4hk4MODh
2+/JuLGbvL11n+Fu6nRZ4ujZQMy2PPM1Xsh1k2HCK6HJyTX05hYrtriM4nkBHmEe
QZtXoPS1pts0Mhh3O34hanLu1BGNlwXwdtKoSTuWen6p1wWvaDuE5tuQISmBgG40
9ZylDeUqVoBN2IuAqo5Lq4WPCksB2660QmILHz9OKOkMMri0P9U64AU9X5Z7ywAt
zOAOmXPGvHBW6Y/NWkZwyDyYEAfXW8iUjmYvW1Yj7+d7fr896O+7bGV72TIWH9dI
5BHIoicEVeBGrjsd4fxS2wltlPIhFTcZYjZn0PF4cumHlP/o0PDE1j/SN5iSB1LG
l5cH74Yq8hnUDD3s1sShCUo5ymuTCM5P854HUImE/iTa4Bn1r/0ySSIdWh2kOuOL
7z1dDiEh063pnQU5KI61j00bec4/jjn1iJGt3ONdZ02H+f9grt3MZteX3gT1sSjF
45HbyV8Cv7NlE8pMfxOv9YHWWqImcgCR3tfk1uyLibvNqU4jm6r8npyU0NJ7T82d
frX9Md7DOysLp156yW4clpyJlpt1Kw0TboUYzJvPMc1lBPA4EQOfB36dM/4o9Fs3
b2thiJ7lDsNQAOrlEO8xvtqKKxYBmCEGcnLLdcVcGNRCJk5KsVngsDOyKLdfoKmt
NniygY4veoAkA11PmaGtKHzojGi+C6uBvPb0w4CjZpDC1BDRAbIqfJtDfDwFJX2U
ulyyX6MGzmS7DnA5MfwT9ofQiJDlc0sbhqYXSoi+3bqYXDrERFILAFcx/sFwsq5X
zDCF0CSrChZho9VWXkN2oVsyyWaOnqfhsktINFMBtKNx6URGcc4PwZKTldYnmm4l
H25E3+p7NiqAUggQoBdCvb8SzrnqWsQNNZGyikBYPfbs8CAHtBevp4xxMc8V8GxD
dmHx64i3hPdRi8/zU7Eu+eMFgzwNL+PK+bpawB8hmRhjmSby/7smaitbBF7W4Eo+
fTe8IRNdcwrUPrCjKxAptjcxVDhSQKNzUxTjMo5f2pucwteB+/SevPxWh2vhNT35
sEDV3qb0YuQkVsJzMbVCcyRKtQcwcuJ6BYSaCizSK6HRqfoEYBTRMNYJPeusUFGm
a7NHwdD1E70ftW848IheC3OYMEMO/BevqF2xo5Vs6Es5wpt5hwOW0g/PjsmSRlCq
wN0tthHtaGTl+2QvA8wyH+ehh78/5OJBBWRKhLPtXMbu3vKACo1JrTrPUaJfW/zM
VuMPxvnOdrHQ+l1HnKKjelUqN45De324Jnkz17PByWjP6cmqNh9saKda8TYgPVOm
2jRHzHGrqKqn9wN2IlI97YyN/HA+myN8mCIbiXGHOB4sw4QdgUOvd7td3OZ+675S
2cIP4NNKqkfdxhOW/SF0ldYUnhTne9KkZwufDe8DqVM75dFTqGozj/73+J1pTTnM
QWceLAx9QBEvnInfv+ghGcQe9G8Lo8YO8ZKElMPLZFfPfcT7xtQ1mnD+PUYcQhEn
WcrOr/ZyRg0LP2sRHNpltDRoVncl4NJKkJ3XcfRrJuTJcJhw6qNrBrS9hSuCKJ/l
tdILZw9UZ2BoGOZNw/pIQFCnLf/Jn7eZIP3GBrFxRWkpXCmKciKtI/IkAAeNRDs7
ukgc00vkmPDCS2WfBGoqUx0yWz7xbSOkNOJ8BAhrHyuXY+uNXkyidQmavuZQdTET
zvk58FDhV+o1SPQawCLMPf7pxtFHn27JXHtcEE8EwitZ3AlG8BThnTkxL9zAYtKC
K3qU/+6p+2wEYbCuN4ggYs31YgR3nvPuHCvC5urBFQmn3Vs6DcOcMHeC4r3yHdyH
1o2GyKExJjnmBtlW8ITcqnWKun6JazVj6+/21EMX/F2AhLqoU4X5dI30sTEqd/Xv
l6tUsezaRcq93v5CXjiAds9lmHyoDQJQf8O5fefKEEEdnASmF49kP6jQy2i2Z4Xh
J21vg9RrVG3pnZUe2UJ3O+eLzSdM4dQ+4KPbGTf/ATrCdSrv8SC8icLXn7tuC0+u
1JwByQ8au3Jrxr8yLFXmwNbBFGy3m7hbG5ROpNZF3Y5zMGAZzjmgtOEKvSwWVt5U
P11zAJ5Ng58uVU8s9HGdhhVGrNF6MXeFUA6dEDTX19NDCDh2TThIsDEVdmK4PQc2
yPvZCpGHJHMqxtLJ2qiOLn8oZY8n99UNIGBDRXxZWNumoOOAocJBKPKc9EINezjR
PgN9jLIJ6pT7jLuhrpXH4JvZC73yx0oUGng+sQF6+OrM39J7ZvuEwsjWsAQdNCAn
B9NNDIj8r88Sm3bZOtWpiw5XrkAcooIST1Jggt3sT3A1LTva3kxY/KHh32hSN64q
FZnhpYPdgva7r0tqszDNITCQG08KJrkxvkyfeuwWC8d/uBgPWc05SRXxpeclDzoG
`pragma protect end_protected
