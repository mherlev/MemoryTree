// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:55 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
D2MHhS8pxMAGfE9GsNRE5Ej8n3meF0Zj+9HadBYlrUPW2NgGZrfKDts5mpYMTp8b
QGvjOqZCHWZGI5GbHhHSogP2ZCt20Xm51nLOoITBTJaysaZn0WQKjdRENNKVioo2
uloe+Hq1WDwxQWZt73jD3UpzjuiTE5dfeJjXLaMdEWQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 46752)
uGh2DZewMboAmxkPQ1Yru8aVFYLvU0Bn7pR8TstKODx6GRF+le7nxxVPNGxTD9Sb
7wbGrG0nDs2tU2p6SPzFLN1p/Bz8bwQSL/lIlgCfjwfKsQMyN3s+SvuB/UOuA9N0
gnivDOsoSpuGQkW+QhV9q1icAIIfwR2g1Tnkxb3wcXO+zhWMTWEl0KdARJJdFbZY
OnSawmEFH++B2KPoJJSK/QsPxeIyGM3Vl9ahQrYV+ZmdmOIjIpz5VJicpkzgI9DP
/fgtr3nvbrZ4gmdcWTQj78AkljrCiSyymsVd2ZOU7fCqV6k/aaxfuZwwEzEN8KTX
Dc1aG0KzNai7aGahagAXls9zUqa6AB+4h0ajgBUrTg06TeBOqR2FCXyUwRgXQlJQ
cCjklAWah+modOPOOrZc9FnsQzTZey92qyKeQynoQJlmf3CHcR/p6Ad9ht/5eN2j
NOV237dHMvnVYAExDZ/4JoZ2iWYzhtUgYF9UivplGMLpwvNeU3Ht28HDY+I9Qiy2
6y6r+Y2gj0PhWhPKpGNgDnh7EcRZ5/NLdq2Mepsl0rVXdPD+lB9i1Z4fdsPqX6T5
dTJcbNvhX0vnCzjyVMM9wndYfwft/8vgQD7y7dkowa9x2lsjw96ZmN7SltgX1zJ+
U2b0oaQoEIWvix9nUiIlIahFN6cdWeEh7HKt4yKj3ITNtIlpEz5yWcfuqe5O4RCV
Kedk7RWiMLgWFb6iUKDim86wWPLyDIYxBO/UIBtxRjyvljCESq/sZG4iIj3f0Gts
fRrHngm1V7d0snLZUrHdx7vYatZNztaWtXP4otVuHkRKXj+brbJOsE90ZBOomeXR
4Fp7WX6HFIhuJXNhc6rpvHTJBjNMgoHj5UVnSGHJUIS9vEzejAXREhqqimEd/VZo
SIr6Xmn/a7GpRHShHhuUfKoxckLKn3jSjbedoagVx/D+V0YBtnjickpMeTzJfOuQ
lbBXkdM/fLDaUYadN4nq3hKn5p84zfm9xhBT/WUTQmOHI2sZiZIYb8i4zR1OPLhG
dij6zrCNm4d3r833kU65pWCQLh/r3earT8TDqQZ3zjYOX/3DKlEVxQnta9cxJXF6
kGwFHd8hp9ZvD35UTc6+tAozRTPtX5HGgZ1CE8l3xWhSUXAI+tSHzIYxCQAZQuAN
UP+MgZzH30/811q6ObDAIhI+Uv9ZSVtdsAjxHyBbe+CVav0PIIIOc9aPBjvgJRd4
g2QMo3XLceuVG9Wq7tqeRjQ5ZK4VumtDqoay0Wkd13LMjiYEFDt1ZxdJ6dUCz4vO
kA3OHuTHLFfNN3cvR7XmUcVhbXpkPEGgWivNZQ6JHxoG2enrz3lMLXjG/oQuVD3B
pHXEYDFolXFgb5kL4g38PeXyvZtIcLawx62thiCFcPDmrCl7VXf/WPYB3m7GxbKf
cLme0gY/AsDXUxAHW4iIsWTuZi/ULU4hur2a9vDvTHlxrMpXCMxcOdyCZ4ZYdztJ
aZkDBsraH+t9Wmg11jnubZ/Uvivt63iuorIWMtiUV/hUo7MK67NG8kdB2zhAk42M
kNhMnPnRfHbXJUKWE7n8LfluYqvuOvBqSZ/QmvoCa4Icih4B4fGCiOrI2cgCXUod
DwAGswX+HZzi2RbFjigrdq0Glkr7mggerjaOlgoIevrjOs0z49K9lMAKleO5ybac
yERKsSR8vhU5dNuEHK2vaHCOtc0MNyvLWg4m1SCSylqdL8QAoyExO+P/piLmP9V5
q+2dQmxVP5FJ0ObfGL/KwI8rQDf2nCcNjyy3SkEOs0xmb+Zu3IKII6KVW2dvhW9V
Xk+A0b6SHIqntQ6CMxf88yybP5XofWDr+TKOQ2HkOe6gGu6CAz94MciVqlDzu7xj
GbdUfBW2qpUBsJrArOImvUKt6c1OgpsDb+NPJU7aZ/sQxCx4p579SAH9N7QtNDG9
T4vyx6WmEjG4FFT6lI2XjRxJ7sMJOoL86OMroi//nRNktg9Doisww8LD/mBHcfSu
j3De+mWgKs60f5+JrEumhPvT/ne/LtF/7Qi1gC/OUMpSowS0fWR3wnJL/dZvOr60
h0AD/UUJAJuFXTQxlyGkUHFkT+gmOvK4IpofVCwbG3hSOkb0p6EkZuaudXv4YZul
8lb2CSZ+2+tPJet4GqogxkTIZinLkv8t6BZBXPFBd4ZzeNDq0w6gjcX7H8fdUXcJ
E2GvS1hsLMCav04fiR2QJdqPJNu9B7ODGhnHN5Or7Eb25atPJ1kdw+DWkYXq0c7f
xjuFh9gXL1lUndUratUz2gK2Gi967HMc4b4e3OASMgQmD1NkhWylo4cv18lBv8cO
/9F+sRyf+fJOo1B8l3chfDtpjP9xCFu6ql3UuOLHHLZ5M3d9MiTkFKVT5SBtLTDB
yrJAekXhhWr60Ygal12ePh9u+g9GG/GwmiW0VUUQHngr26wkrhTgN9sftp9IifH5
UBpmmr8GqRyytrZFc63BtSRDwZJm2JZnlJSon8GjVwexPW6wTWs5k6+1P850nT8v
ouW32kt+gMDR57pc4kp1RTENi12gDMGfQGbgAj14WrQCm/FbRnxtRuDbwFcaNCfb
qYR9hM2L0HytsUwr21tgm95lJ7MMrI2BgnYAKuUa/c4UjmIJe6Q0+TDE5xHrnz9Y
s3Kyfq254JwlIK4xa7mCrlCiIdyTX9X5xvMbd1/4dDc4X/bBGkzevewO7GzP1Vuj
DEjKtbPvyRvGmjXPf/MrFTgvZtPAnvstnbGU5HbWKC1EWqWXd1cpJccXVitCvKmy
yxeMKVgeEi4OGc6LoxhzKEhM9DPWgU1omEqPZPaybgZm8W1Y9QMcaysQ3fJOleos
kjD4wSFLVZfgCLKzSrxyacHGwsP27HgASzkAV0hAI5P2ZWfycLW4y6kzZJaYC9Xy
QFPrXVk0DSgA/pVxZQHCHVI6pnn0iic3QHpohKdsLCPB8eGn+2R08cEHb6Onv4X5
7Ik1fa+F8LM+aFBJF04yZnpTru+GzPzOlanvpH3Ja2WumfYvze5YqynxVU98Pr35
Ykwz3X7ZwGKae2YLYIjIo8J4o7Ib9lM0PwCY18VHpG1g36+hFFDemwMDupRaSOSm
w0S61T4XF1PJk8SI6A3TYFfH5rI9Z2jEdnUdIMzGOwn7KFYTtspHiJHdx5d1FOKx
u6V71K1YkgCJVcFKwO8o9JLdqb0Z5hyCb9AqxqvOp3hl4qNcCR+ZQLiR7mXqqD9e
kfaUKcoPK76KpLnUkLSus+USOLdOk89a8uiBE7u12wtdf+5sD/cqKwNE7uiLYA0v
kDTvqx3YRyLkvXrxmSat2nhKB3tQ1tFOIuCrsZ94VwIYtewdE61ExvH7m4uZJ6yj
D9sa/0IrYab+gt683Wi+Q+xryDHbML7qcD6ulKeLQipbe8F0lpTE2gP9dI1f86oJ
5i4jwJ8feOvoyVFn5jaSoCphDwlMdqbB4VzODWEqqknPVNhewkN0AqErHGnyIneB
ziEfS+KZCCigLkjwTbJiyVEt+SQH5Q/D4kkNBhXLfRoTb7iSiota2HxSJJSmYloV
Wyr/+lqqCW9rzXdT4eE2HLiQb/HvR9e2tnyj031URUyy3LTazWh6ykQQ8TdpXZSi
QDghSG38RC7S1BIsD8IdXDhKOPpOJf7MNQ/b3uaHu+62uRFBmVLS6iTY3Q55FCAs
svyu//wC8WnzJwb5QMn+HHYBU+Cy+mSndJM/YaITe+fy1yYqOVrrtL7v+x5BS5mn
um9FfJ30pDjB41JW6JgBJLaW5aSziSFeGQGnHXCGY5NOv1O3wzTiOB7qsDKpOQ6s
eNmOQTw+Hum9nJ5svAXyxTRRgFnZ1I1BXny7lOHwdvju9M2y6gMkRIdXAdvsFnHH
G3pwVTjQGutjEkX2dkoGueHraB5WKZPUYPDeLrm0cs0nXb5CrJ36my/8tLxLvQWe
TlGjudeWINNcwARmluRWDQ3S6oU/NxnkOfYSFfbdr+FkS75gQV/hRc5Vi9x3ycVj
82HAEuHR0KtxZDrGxLW+2wWhBy+0mLBt+M6GK2VTWr25zr86XMhU5oUtvjYgrP7v
fxXYzSCkQABR3Luk87wT7YM6fSb2RVioxP6dzin8z++4X1zzBJsYBPH1LzqpOBmw
qB6/QqroeoiWNx/3sbvg3SFJxkPRsdPHDFZ3EZG2FcQKKEw/+E620xOFfPtpvf/e
JIk2uj/vcIjkJyAZhZyC2TFMIN7+xdpALwuRwwLOFRma/m/fxHD269PLWPvNcWtE
lkUF9kqply0b0DJbBhtvnl69LU1nAUWj6iJnJGGsxC0pwClQwhgnPQ8jcdwtBRaD
TdPyDdz1guTVfRKV1HlrgdP4YY3/UMEgbr7hgMmca9+LIo/C013C/8R9IW9av7Hd
GLW/BTPKZHMCriBT/2bF5mOsw2mADH7aJkEg7g0ZIUhRfiCwxSFtKRIiSpX8nXwQ
1IpmweHlrRXoOdvMS6ykwbUtXJ29MrHGH8Xeyo9pnlcB77764gS5EBPZzJDekCHJ
Uo1LmESMpkHDxh2YLT6KTf+/PfuUMOODG/sP1f9+dC4z4n/8Y+b+qlY6hDS/1SjA
oGdVH1I7FhIA/NCCn2THRA1L1o7S47u8dEHkhLGDUNIULPDQtZh3ZJh0vlcHCq1s
kRhnG6jk26/M2W47utP+HcP6M2IcoeadLaxYdTk+aSMGB0byz8ycaCI+Wz5PlrEg
KfIcXznAdo8mMGFq6IFMleaGFPQK2bmPS3wGSFEojFTqeHelzBRW7IUfT92AukcK
ase6S+6vFL2DdY6aVkMH8MkMfNypDj+kZrJAXVRajpdtbpoRDFYWeR3QfaGKPO5h
iJAwl+7mvVOXHBnG265p4wetwFZJNLtDD/BSe4yI31hqoqKyZ4085P5+G9HAss+3
pnUt37MAMNJXJYFfJOc58VI7mwi2klBtCCmuryTQ76AWAVq85EoESnB3y1wzapO9
qCZ/IhdnW0DMIXjBpfNJz8Gc4k1HV606EDbxD+JnCp+x9uYWboTwJ8IE4Q8vP0m6
U87DgeHbGMTB9AhOzlv4+5J97vLG+2DItZGLx3bqo+CM7rPPQLCjPPhfxXKe6s1m
mJvInCUcjZpS4okYK9rNR29JE7bkUQO5oN3M4kgduAO99BqC7WYud4dtEZqLF1Vi
TFcLPNVqs1U+mpYWTQwiJYhDK958PKvrYdOa5cUFo/GyvUFIQsRY4MLqJ/KqzGHh
dwxbPINjAU8buuVRFAkvcP2ywFqb9sYzQ6T2W3g65jZbf4s8MGDdj7GCoxChVspc
jd+VVw7ZctbDC41T0xWFMJPPkoYhr2YR2kdIOm47lsUal/Mj3A8lqpCMLh0KTI5V
LZsMlCBRBvZ0EAB2ajP6A9jlTmkdEXB+3WAe+YJEOcXqiMSPUp6kLu3T7BMneBml
21Snjd79WL+zEEqjBYHXr38laFO/Xu2PJPp2+LtXpbi3tqJR60TF5f5VIYU9a/VM
/o4fp0e7W+05uh+RfM/RNU37qV5QF2eHEiZbYRnEWtsqwDPSCWmIytnUN9WzTrXV
oXZbKSHmdOQs+HA7ehPHPdK0DShJDOlm45ahU/vjjdTeHLAskZwvvAtslSh+OITT
BRx38J1iRlu7xMWd9a2W1CDmqg5fFDkaN/ylTm38THeXoFJYB34CmImiXQWgw+qo
/oQO4Wpfcrc0O9GXdH7whSFuNPxR2S5FUBQI+9IlyTg8LpEAMMoDwdI0GEJ3ZrtH
+2ut/amuUoaGK5Ar187TB/WOi9xAQVy9gT6FW2ArWqAA4KOLfU6ZgRoe0LbYpf0y
G8LyyU2U5VvYejCWezz2fFCXjsYG8Da9XmLTB++wHj/ZyLskWQMKflIus3unKiUt
goLW9kWnDOMHuN40TjGKZ6WELSbQJg5OmdlYj8LIg7IYFxXWxIiUN4lH56kppw1C
bt7StyHhQd0Md0zYd09i84OT9nAh6NiwgZfZv/ZB9RoJmA9PpFdisRFlnSDxcIKr
HYiQdGeEGT/qMEUJGvAhV9uCqraPTKyBjt0zsf4V57DSB+xpesKnDS6oYZv3Z/tj
LH5RnA/GdWF7crnhttfPK4DOkoQwK3aVpDsjLFwmoOk2Q5rbmUu8wgurYeMwUlKU
4/10dOSjfQnfixce/rq6hsjdBlNfbTlYGsFyW6+oJKf5ZzLQ/E5jw1J4rsJcVBsR
j1VTJ1qON9yqCT/QESDuwin0N1S/Rg2Cuok3PRYdkTqAQX9EugeDn8NfbB4QQlFN
CobAglkfCGZ7R6jWyKuuxDL4PEHCl1FsQF1BaYD7VxCwAIiTwYXwxh6yr9rYS4dN
CSbGTwQ1p+41dFD5hwPtTFLFAntfjqugUs7VMdrsfbGOoeuTA2AQpFJIrHUf+NQ5
iYFqFxrfOLOSH8nwdYpRemqnUEFwjbuMREuLn+C4fKJTyHiG36Ty9heeI9SAu0f0
6oAyBKQ48uhWaAdGUlkea7Vxe8WgaWsMoiM4uRbuQzw0XHS38j8xr7s884Z5lvdX
/bpSDIt7hqYi3QmUGvXcNxkjwu9+/tRGjh35KnM8PVe0CtURZDqAPxKhkRY6n2HN
FEv4kP7CRNW6jTzK8xjSSV6rA/0+Y5kg5tvNqrtn79nNQcPqj/mZKMwwe5M0ShQq
Pk3ShxoC801mc+212k4jBHLt29HkCaKU8GNwkvOUY3PqiYPLVc5C0gWUjlYA7v3R
AkI9iTuVOkLoWMOQeAsCP6gRbKjpN1ExWDw/IQyLpkuhze0UaE2ZVFjEelPwZdP2
LcWI9w0QeBHLdLG0xPuihcqHevuSGxPtBR4ynKldHIXVr3qWq1xvUxrnuyxqhu9L
kKJuJshvPejTdDj16QTy+NV7nSZAkK+DsYZsiX0OJk8wUarAdRrGBrMXS481rynk
CtUAftd3APO3l3Z3JV87GN//nEJiUmc+8aAAyIgYyXwVxVIaBDJxNx6G0QPkXdMe
NcSWymQvhCg7VT0Epg/ItHNi+l1FSHOB/6kJZZ54ALTd2nkEZsOxcaRD+sDzgfcQ
v6QkCn4b5hFYolD8R2lk2qgh6mIpOj9H11VqPU/YyFu4ZR6hBYEXvl3C8CioE3nD
RTjnGQT4DHZwkoQVkuIC5pgGYa9JFA4wHnVhj4yD94Cdjdamj4fRxBDEIH4KOH3l
bOF9NQZ1sC4g1CfqpRPx4aYrkyTs70SYINTeM0lt+XLzL8bQ9sU+/aQ+mYCcj9mG
HdpRcNKNqx3RpD5hqJ6Or34bYlKcidmqWQ2pc+A6OZra+A0PfB+JNH9gLZrsxBMa
tSHEtFT7u4PSYj8/okRU35/zyYSWLrexsp87bGOHeMg+stNNXjI49NYXMLdwO3oc
a+4ADaI2SvQZRByaR4XTvw/BAKKB7sfV5+sVMnv5TfuDCRBYLSCo2Dv28asAdy1U
9NERw5myaJyH1LmivR2DM5cN1/Q5eOC2Ngzrs4B2oAOiqf8bKAnEufXeJ/Rs90ph
UP8MKpML4ZLN7s9WqIc+r3x8en9fJbRONryi2UN9+nsvDuD8Xw5c4coyY+LfFZR+
K3OTplce9Lc6ZdWGu3dQ2/tfwRjQo/1Mf2zbq8pvtClvwO0X9UjcjrmLalh8tGeB
vIQmRx6iVUyH41thAxCSDmALWRp5jXNF2o2Qg9gxk07Xph2o+yNZMEahIio/809F
ZaOs8AePG3o74QxIorkhcSHeEpgSPWUsRQvxgArRCfnd9gLvQOaV0YC1qntY1sx1
coGx2QHOSI1eihb4chzbUvdRkmcCQdvVTDN3BU5vGnmhTxPHAOLcD9MJSuXZCOo4
Dfog/ma9gMDEq4ZrVBiOU0SliCv6s6q4ky+JMAsY5pNqfCXZNZWEgPm2Pe2YH2R0
aUz1gn0dzvutzMySnEEAcGepP8lx5FePytqsQXqKDNECAoTbfmmONspHxD4XIGgD
2pTQ5tJnq7L7nOwU3xcYKJjsA3yPD45jPF3yBYZhV9ZQ2PkwJ2cxNnDvCJXL/RCl
DTSCFUeZEJxk/l8nf0vjhhwLtPXorD6pLXkoIidEq0UJ9P0bf0YizglfFFr3D1Ez
M/KJtlpHl4SrkhREr2MD9vSneQnhSFLt49Ntlre23UzIUV7WCvbn2QSR1DWR8QpU
IMgMGHE1n6ZfY6veac3UJza/eHjlwmnVfsPEqxNLLWp76Vwei3/pjdgivVnWkYn2
J3IrZnQPMG2qyp6Bbw059DJYlz2ETTdeDpeFUtfnpIVPxqRftM1xmNsJjCL82Sku
Lqj//1AJnCfTRO5qJtYH2xeDT27VXiQ6NT2ntzddEh0ZFH0rwgxXlM6TU54UJhx4
v6hgrwufQCEo7zd4Q7QUXH5SNgEE1KLklZ5XxJa0WToDh+j0Iyw1kSEvKk5NPWtf
pgBuqU2N8JIE79/FfCReDnfwzpcPU+0S17AXq3G58gcPUx6L0FOA1+qzI9u+6avq
TRQUar4kUmjh+aXa5bonGSO49HOVun6rtrFc89vWtgOddqqthwUBWOa06FhvNoF0
jIi0nYo7Myz2P5B6yBg7IS7CLnkktyrw370oOn1TYOnA7zJ73uIgrKDRqpGcIhAW
ihalboCHf5W5d4s08PCDkypDpPFRbrod0hNfDlQE2ZAKYcV6dxywvOb1lE961jY8
fJh6vGRg+gQhCWRz702HgzVDCmpHf3z0DtnblFYpGcr+YBN0HyIEc6AGceo1NCoX
T+RENR1kJcevzEDPtIq1XRMC9X9812S9JoTEz6aNTh7d5zivpSXxXmB+ICqKNNZL
4icFMF8+2aWOmDF5etdu835sl75nFQyQi7vLMy/HFm1xUsNO+skYcnDgOwRcNOE/
LblkGC988vSCTVeQaI1m5PzPY84ehHFpKsyECakia40gzjKHGBcgTQb5hqfhNoxP
FSuKP+DJEWK6QGRtWXTCOWf8VMsqHGSoJiww1yGR4kmDYc+7uxXZfot9FGvL6zPe
y0e1R2bumSYJknbxbShCFO6EwX21/z+qdo7jco3Bnrau47MhVgfwngt/KUU7hhEN
j78+GUhjjnPC4f61WDLSju69fE8VdsfntJ3TMM1jzliekMgXta+RU6qU30aeRgj5
+M2t38d72yalyJYERDHeGAb2Z5jZJs9KE7mrxAobSCR/SmNByiBNG3KnLoRIOHFB
+5bXCdVSLqFcsu5OyGWhpAgHNdarV6MeTuXtjngyAZQUpKZwbDqPPxaTx8wHjav1
2k1VJ7DlBzZLg4rUcNuNo+uHjkvRL+BgIjBgN9faDSPbpE+IEDjkoTgR6pZVxnD7
/gznqpKBKmzeq6+vbNllYTzS9K/q9ticCErk/tLlWt4hRsFHkbXuH98qaTWZEfx2
vHQwj5iWIweO0HcwEcDADizCOEXP5OZ0PBGBuwvwEsb96F1d7mkQ2nDBmREGVEUr
qk0+pWhiVyM4Zku5RS5Q3MA4/y3F8p8Ywt9BfmNXbWM3lAtcFV9cDcwl9scIeZZz
gtZEvFoQbjWHMdbnhEsdeDoFFmNQJBJ3r3Rk44H2t0bgwkeRhMzTS4zksFLAyt/5
siJC2KYIS0takWHDyga5TMzgiUXJJFb801ysWKaM9ly/V2/F1BvZ6Xj4QXap0n0/
zv0t5n6QEyHvpe1EDgQ4Npg8PKlhdLQxthvelkJuEvQ2++v93BAnNCXqoKBrk2HL
Tf/y/HBlTI2P6JhvfSvdX9q/ReEHD+jZ7vAFzk7o+3jCLrFWiFdpsJF4U9FlJs+O
VvS56pLHKH7eutnKSQK46OZvTxl+ef6eCPhx7rl6ML7kBvm5wbEPT5Js4VtX4XD5
hRbo+RUHX6cTcy1oQkffA/dMAN5UVYLf9W5Sm8+XIDFwW0KEed7jwLCNzRr22xF5
hmjN2H28JZv0c9WwDLPMAVepedIypm0ixdrqfrHrh3jf33RA5JylAVXO6IbBZPUr
IRslAVy9DNVH/SI7RSEcuxmvZU2il6c0nHNyR1EzjTpxBVsSZW5KPyAFmAmhkNbG
/6/mX/dkCuQ0/aBiSsGd9hQZdjef+k8vrQu7a3qJO25wREyUyEfeBK4cMqN8yHbu
3fA/2wudqUE81qbAY0daCKg1vu+JqRD85VJTeeZuPHVFnMxG88kzoZ/UC1PVnChU
c/CpuNfGjrnd85Iyi+a3v0gGO1w8JEDWGknTw08zYBtIdgOVOzBndqLVA9+BQpRU
y/ph6w/oTIqTK/mhk1iYiTF4us7HC4BYh9yaRbLQhFo+nU56FiZ1jrb7+CE71fKs
eOvIbeuV6VGEGpE1IW9KtSq1gfvahQ7aKGt7kz3olijy30pkAYEltVyA2QHAr6R/
g0Lpk3mWd9fa5uQnwCnszJIZ2Y+hObJvfcRN3b1wn0k08XIZfntpL99LLRt3AEuY
sNSUitj1CIg9RycBdSG/nJC0+QK6Fx7uRrq6FpxZwQTDHd3Tc2+owPEI80ipyJYj
q7s6Zn1lS/z4oV4WlDhquUVM1gVfwJ/yIiYp9XAMYToNIeyb1HWqa41uffiEOlGn
ih1RvHb28JvrWap1ghPR7muiXXB6VQkd83gSX6FxdzT0Uc0iUltdsQdjdOhJj0At
dL01Kujj0sWDbppbB11NOzYNl1IM9Gl8yHsGJv1Wxca2aL4i1yGt28ddiN5W9s/Q
gt8qxRcsJsPLDUFLGaSyWbXeOpBEkvYiexGJSXnGIoUldgZqgPIwhteNYAnym5m9
vQD0wrDpB86zeAnRZaYrW/jCumbf5G8uz2csOdrHQSzawTWZTjuA0TV5jv4oFvRd
hsT3wHTRRVuKfgZK2/RzpQrXqI5g9jhUIBwwQBqXUoJCGfRVA0Y2VxgtkQfaiWU5
IIsgE0/hWnrcj2aFkzL/2fjbtXkQTCwX/qlwhbLiokXyeNE5BUUixmUw/IuKHFw1
9Q29DBx075bWmbUrSZrAtxc2q79qq3UdsjRNMjmWxQpIbI1OaQsaiFRk5oHeSael
sejQejhiLL3SeY3mhN+Dq44uW9hcR1IlqKs1xAgC9+64LIemZ0is3c0o52X0x8IK
xD2IqPgnI6lZYACvQQd4z8kUGqbnKeG2YxbB6WxBtA7O+MxFxeNhPiEj74x3mvoH
aH3oxqHgLzRbjxrD9AH5Aufdr2dcmKVJou2XdxM0WOmSGnhUyFjwF4p0hQmUtDEK
yi8TJYJQYO2F69eN4n28XiJ2nOx2w/Ziw7KShxTyxB5/Au88+1IqMBl+UWxW5+vD
9+27jvbkHFwVBm+LepXe0vhrtbYsgePxH0yC1mmtQ48jNVFsCE7H+L069sPmUe6s
DDM9n595RihHwHfUzcQNuejuUK+9+mHKvuGFINbuOC9D0j0f5PViSxeyYgFAhxOw
gDkGkeh8+AAkJKeV003bKb/YCNX5OOwWVSC4yHualWuhZ17KqoqabNBi7HBKDtxX
JTUhs15Kmeg6zh76XuolDzqUS/9IQicdSL0YnSp9zkrRL/9m00OkQm8SZADhBoN6
LFI8mRopDjp6BtWxy5afZjWnqCyw57+t4XGFc6K1UlSv1EdjDwHR+nEy5UGgIvxv
kL9mmGexFy35kFCYUsYpnflQoUd7Q+aEl4xqVjdllVaI92K1UY8SenZaZZtBiAsn
c4geW0PV1b0wSXbe8QMROx4nszIU01jU6bjJOfulZEekzNtpEj1TBDd9OIeAV9ep
qSTKwUdMXjVWRZI7FimTOIN8w48cH+ab0K7kxBEMNc0tJBQ4xgDeZ5VGS3MwaLJA
4m+6YnwyiqoIR9U/OIzfXfVTm8By0R0WeJQjwT0aSga8M4p74HGtNo3ciGSFe1uN
EdDzGakilMISYQf1nQ60DTCdSwFEKdUktr9AzqQwWj2j5QLdwNFAmilW42cAcyAu
fUjrFqh8XTBx5Orq2IRMq94eywTcgYwvOtbU6BLXi19ntaeyPZVyU1j/1ZSu/iBC
41xtk/cwK1/0ZpUYAvXsRESCqL0jq5boW6a0l8V7coeZIDBUAYdRTuvk+vORVTdI
GHCTUarqAE0a/pMu9266lZ7cu7PV55Cu/BvSNkzPMOl9i6A6LUnyrmK5A2TOyNk2
jQagbQ6SznkxoJ0MP+1YyIbXR2WiYs0v45MLk04Zon7JI/5tYfhmpf34e3zcmijg
4h8xfSkQBP5TXlwMLEwThrwBQm3fH4lEvWGAivAZfHUORg85G9QQLXqgnVfi7buT
MiZMwj56fJufi0P8r8VBf/3l6cDzJEOBXanFSmdytMaRAne+n5YM7JWHZsTcT6/r
pEUm6YRAVImgiDMeG5e3zELDSgku/qgoYr7/HX3JGiFAryiNy7ZsD+ise7p7Hbpd
l6V1lviiBXV9Z/8jV+RiNwvfFtyxApIzCEbtBcUKYeY3DE50bONIcQQcJRd2/POs
ieDJ9QEsYXdBT5GmAniyHBNQVomkfztEUyN+VMO6s0APqvKKt/3miSmSh3aZzsRx
OuMrli5A2Sb0yVKY0cMcbOmMMjq1Ppg6uJuPb/Tf6i/pQLIZsXEq6f9CBNzWQPT1
ZfDu/n8IDaLBsN4MxJl/rkHYiNoVtZYWuBjMk0U8hYQezbakD2uTsalwvcEPVicV
gqBchRT0MHXPD4tLySBD2Y3911QiMKS3KKOAUgJkRxXUcyV2uKCB76KMmTpZTZOk
nVMclq8wNWC5digFCEDpWmNBP+rOpG+sQSgXXyyXGzpdvprt8TBd88/1naDTn/+8
LeHnpib0je7KykLg/qhbiRu+jWA7NuHbizWZv8Knar/WtU6zITHbrpqCG01MbzbO
2Chsm4CXaM40WcHR0/LDXiNXXrwsNoJcne+2/W1jMN6rjmxfcSrZtt3Z58Jz8iYi
BYWSV2Jd4OKuC8o2f+PLNvrokJ6wKBJNOYUmRauNInx61QHJ2utJobv6D4QQE95d
FiHQ1tKDqRg63a62TED4Z/nzBJ7G8KUn8ooLlgOLyjN3le96RCTC3oshWHcPf9uO
F/M4Rgw9Na/UWE1vo8U2xQnRRNPVspLasXTocfHpx5g3I79YCSf0gx556EBoweWV
1b4314S4o7O1A9Bb/hB8QO+3xpimsqdhvfugBX12EzvM3sGP3ineZBOn4k+XIEkB
CcCo+uo5t4wQYMtegObsRbjrEewKtLPHpD5Vj8CxJ2j4JmVaarcp8zTf602NDQ3J
0ElXI0zRqowwPqPHddptVR9XDLmRRSc64Az1Y7sWToU3KUjTJJnUgdCsgbW+fly3
GJBtfj0Xp7UimugGcQWlpbFqy4UB9MOyJriwxhySSwQ5tAzG8m+xw+i8hientDuo
2FgbZFxYNROaBOPRVP/0q54q2zdLQoQhEYe+R9gjV+nMoJ6OIEJvGhTzLgkjO71U
WRam+u7zenAroO0aHrVUpOpfEFMh7GcKQx7B6a/C/wGin6G2boakVp/5VW3Q3yKg
E1JxBmFVna4CFv5hhdy92Fn5WDZs3yNQYHW9HnBz8GM448Q4K2Fh6bCe0DnEasU/
12+7zq39ILxdebuCLTtZCuFOVlxWCiPExbteB7yKMmHbyfurJKsLVoc3FjPjgkzK
kzF6TRDxNtQeaqez1Y4F8Qb324gvpIuHprM9X2djiwAyYXC1ZREBlrVOKMe/guji
ZZgXHn3BU/ohQm+AqWLgFehvkdLrIdBxdr1Ag4YpN+RyMjKdP3VgvNtH7mtczNTe
dMxFP1g5DByJuxSQLba0n6QecNoEHzt3znDxWnm9I6GOaLoGeoPh1IjLcOmjkWpv
buuHC1rqe4Skul7+U1E42I8j/4F3zUw0yWYx5HLateNQtyr0ghIRVHKMPiAD9iP8
WN2VnPyEgl3A4/JW5GmMrsEMpuQqiy4fIeuNK6s46ji7hhCvubJibwucM97VXO+r
WRfOVM541/WLGS2UDsGNAXXTNODYO7/8UZAj6FQrfxNnseQuLxJOFgWAtHXGHsZV
oXZrwgcxqtzUBiElEexm82tquyVrzmu6hizUHUp0gdbZR2OTNY/5PkjVfjcr5C3U
XuSfXOQVCa1SkLuUJTKQTntn6ml2DbawYJpsJgVhmLgayiAL6tSL8KoBcuEFpwK/
ZORBHPg3TAzBzn1+2Zo0UraEBlx+ZRGQs3ldjDr9EOcaIq5bfr9qjxisweFULygJ
dSQL9gKiDFUOC4aoMkEsz2NUDlSVf9hJa8PxvDDM9F0Rh7bwtqjSRYmvM6pMx8IP
/pjQHj7OSqb1VwHVIPR9/mdqT8PXnaVSv0C+rr7WJn8Z//Ql+0inGiQhXoMOfo9O
pbkw3Gyz+NjB2zOAgXApAd/j0aHbSO15rXYgNLsUYpvHhCemqfcVT2cJ0U5G0aPf
IfSVJ+6fLFkD3aTJWHLQF/GRyZ9SLhBt/xZJ9cn7SNwFoD92CIE4Hgb+EtBgQ9ny
82jq+spDlECVFC8Nl+gKzKbzMi83+dPG7bdSYODVWMN2f+oOennZ/igM5nArOyHi
ra5EGlS13MW78CLkKzUxWKPrUcSPpsD766Lb9hktZjA6S9CM3gSOleifQu3qyu8g
uGeeNx5U/cXWMe6dB8Ff/dcnm9rFWJClDW5B2nDj3O8OXnNBPMjAF/I9GMLx4vtz
gAJYhBdKzi5+fsmv+fNQ5qPa3m1hk+8ztBrbG6rdQkKZCRkMUaATatJ00MMhfnIK
p45b9H+efpwf94geE+dA8ovguhA8NHRl1xD3kXgSZ4pTInT0ou/jDh28j0+HHXBn
EP9iKVi8Pw2Pemiv88ER82jBf4PytNexAUjXmr7dPrrj18yKLhg/xdgTl+0bUEnq
yj1v9Tb2q8haDHjSVqcgcVH6DRuXpPZXEKNlvGuncBnzmaFYBjpSdWIkt04rjcAp
U9J2Xl97TyNryRXAbTPGnEKbgQAyHRsgreGI2zM6RoWtWEX3/f22gHvKhruOdj8I
VGQ/MDwYW8i3fNWv9W7nCCij/v+ojiXqm03E1W/l1M0qP3x3IlcUpyRrdIvsYdFK
ikifPF3OJJyniLUdPD9ytsMg9hEeDNeRfTT6r1LpesxSZe0cx72AJsu/rALGaAAF
Eobw3+waFosyF2f7tkCxMQXgDHBwcSmy1r4lo927K6QAjdo6y6aWNxyrhF3g5d34
Fzaqequz57IGlWJH4nqm7onODeqRb+sDudNzeh/ICg3/MEbIiqZ05I0sQo3MCxcr
UaqLROzZOSPc6UJJ69G1JtJKWiz/2sfEXM79/GTDDF8tLtk3YcQOa7b9p4iVUm1k
ghieggmDFTc8FBO3gFePjpRu+QE0+0Def2JB1vgBQdAVxy84ZO2/jVGD0hcg/IvC
QdLKGZigENDepS3DzI6Ce7NIXkfOwiEu97Dnhfn6lvauNdMyXN5hZZIG1i9Ondgk
3MvCxcqA7lkeiUflVGXqCU9TIjt1HVFqa27R60F3Ae917RbMPQaZr6NDYAkyE+qy
AQL1hIsAKelxds10zeI6TgH81v2hKzWwMOpqp5m1ugF8EYEBGfLtuLCD1cxbdKAW
4wNjPPxlwgSuOITr7iI4KQ1amqDFo8tSmQNgvb9s//xJNsKeG8NAhsnw/VQ9HtX0
94PObn6XY0FZrxZjqBmAu2NIp4xLDqFER4ylKCpojn8uxpRlLaateE+pgt+pMsHU
W06Yk4yjAeDz15o9CfqZAIEtQWO9xFqi6aoRIu+RxxU3BWR2U0rkOgcuumONAbeG
5SsbaZOKGLEfJ5ijU7x3alfdbQAZ0lISW8nGhOzRE2ChgCnUx7riGHOHmgIU6Gwu
qPRJZGlnlW6mm60LEWKVnUM9DmGrE4pmRbJGch4VZTNDZwE11TgslR2MUHHWBCCT
8z3MK4ZiIvu+nwcdUAddrPLz2M7oTFoAjGnBdS8cSfyYZTYEDcLA3xfVMA1IyNN4
QWFhO6Z+RqV7sXuhx/y8KEoRorfNgA/PGc3P8TEDfslq+MyClPJPRSuqwagBrRuR
zAi86P+Q8Q0mOhcQxHGynMiNUiAva5bStAY1REkz3fFfuQEskbrCVIKPvXY9ua1U
KS/WzMsqFjBRkQaLOa8gI+mh/ASpzKFs90cEEcAC4qCzcj4y1pBKrNY5bl45s7Dj
TN7QpBxrBwpZYRrLecjjBkw4MbDn2vY3HxbssMnfGHwN5nx74pDjUGNnl66IaF+V
8X8Sjza5GrDgItvw7tr1GkXyXN9vdB/+bCJBT0fBk76oHcX/1My1nVRMyOaxBktJ
uSKcSfriBbOhix3dYVHPy6ZbNUAX3R+duA+W7rpSUFf/JgxmxbYWEDfClrgVlGFu
F9oJHB/Q3mLoUUK5IBmbKWu/AZKL+Ejx28pLY2ARiEHtrTwFGlQA+/i5f6VmOetH
3xSVc+fGHK/8I1H3ZBNXMgCDT5O/z3mIFLCDqbS6yAQyfmEUVPBDJrxwjmRD0mpo
wcjkiUtuY2gvqDbuLf+5X6r4cmu2EdbIKiDUYG/Tjsbq+HH87fDkIERuktaBePvy
8LT7NbvxZe+zKJN2teMSBk4OhxE7K2ucX8pM61gd9czB2p0YVLUn1ueO4KuJdvFI
h6eYIYrS/EuA/YUWxLIH/hMA0tfCuwI491GmbBsEpfNsUzbXGy6vxQY1yWErv2Ej
Kl4L2QnnmHr1/rPECJ8DImkhrhJSK0PwlefHblWCnxEVTtkYhASujzf4fofDVlT4
SGAbtLXNcAsiM9E//GlIG/In0xS9f5bwOH9uQfKRelCPGmcCCR0j+UMyB+53qoLK
tWZ+5UMTQYp+D9CV4hJ9d1jwWtdGGQ54mTUhIGuCNvBxi6+Nwx09Ijh6cW68Gcpf
PH158YcsoHNAhjztNLSYEl9MnicW3Y9v7VooS1wW682SqLTOvkYo6L96BLYELo3J
9KvoWL6uR2575kpVcFQ+3Ko7wmzN97MrWlsR834+ft1ous5PQ0dZY6E1fY/IXkTe
IS3IlCbcwSYMlLHIWec8vTb8oG9Al/3Vxk01Mrm5qdgTnfZ6d8ZtUBtZ8BwejV1p
EBocFW9JpIKr1C4ERyOlAR7MPoOQusdZ3XQ6FpdFzncBYj/oykOAHLKCYJi4mYW6
81fgRZUJIPIbGVMoBJB8eNxONkwuBhXjUH1yEL8o6wzYp78bNQ88SeaOqJwvYl/M
oo4jKuA2MS3Wz1QOeHsgQczFxeFNspulSyvaEpUsO3b42deBXFctONUYO5Te140j
qr2ncyv+MCR4OnYyo99wyVcnOjOZ00NfEHg9vsN7rHuMkxnC0c0fd7k0KD0G/Sh1
DHQlBxwyyc31ERA3GV3EVgWTZkg97tieadan9sVISGlu4zn/7j0aQsVfCmdWVCM1
9J71TjWzuftjvNpwXogcTCQ0y6ITgvWenHTDw0kSb4mVwE67mBzN9Q2IGzpkuZir
0y+9zhC+6lVKMwuImT2IYAy+ocLP6h9E4w2tIs/jZ0w9xC12XQchKNATLsNIjRtv
Q4vF4ois0yMxGOyTIMP+5e2TZeDOl2rCrdLUwjkcuBq0MYOcd8BOsn6rU8xlTiX1
a3F33OmxhSM1uvb99xzbnWLfDp3CasOXZ6YHTDgKG/hpQDlD2DT8aFfsfdKPYzDS
ha3imzF0Lq1U6hEt1A2S8O55hJpWPLHXSOWuL/MeAD5BFcZcC0qtqwb8mmqNyzZJ
HJtVtvhx0CHg56lyCy2SnJioqrYEyDASvBmlZjsbXPwipwXNDs5mlEB9YszG/iAh
WeqwAyLWG+aow6sV4slWnQAnucjBs53t1VKa9U6vTBw8WMGBaOfWxdwpBksBL/h2
zjIr3AYeQ0i1Obbw4V8sPR9eU9nHcXufyHsRnmqokxiFROqI0H5xpYJHdGVeKYxk
twN/cdZMQFoyEq4WSAStaB75uusIUSFWl4to/PQPGn5FNTBZefB0JNewP324MaWC
M11LRR/l/7IQIwRcIlIjfjvx/3EFLnj2dlFpCKgjr3Lsl2Q9W+ioUB2IKs9DEUFQ
Etvm0utKat+BE0sJHsolYavdjPalELYc9i6zCj2cfVfCS0mgzIav/hMuKt5Rl01t
K7JmT+aeOlEBAPSPBj2377yhNKc3HqacQn/UdIXOnuQ7/nzwimRAhsOEMmuAy9jn
WBmaV10kAI8xhMlh1+r6pPMwMtT0iGg/oXiOCC/n+6kzLUTgTYlittidec34lD05
c2KYsvVXFDXBdPORbm0TO3hOLSdQm7sG9Ctdf7XJd6jg0+fwT4G8o77iXeGxiSv2
Fu8vZ635Xu6SbYJxHPZ47Rq0eQZtuw2f2BBYwDSlNA/4EVxHZpKSG9ThO0rq0suH
v0lB8VGsXj+wK0ZOJfDnaL7dshAgyceInxAEAAHZI/6rCC5MB3z50gjwyg+VB0P5
HH/GlMcywy7JpQiQ0agqFWnYDB6E7KdY72eiltW+iZ9QZyqFSqBARRL8xxCjnfam
F0t93PNyhNMKBoCTUlUwm/fPZJcS8VtKmaY7lA/xhKio9O1UpdRYeICZCY0sPKtl
y+xm1MDsfy3+HzODuGz4RpixNSt5/BCLujlZoBf7tfKabA7+LbObfRot2ZjEkpiV
+sAzvNezfbRZ5FH0xeIkoMS7kusrCgy8GyOoWDwB+G/34Boz0fNVJacqHQpYPrMv
Ntiyahabv/0VpHD+deCImUnWKe3gAcXZ/cfMk7PoFjGrKBo7FxjyskCpg9iQEPye
gdToiN2AY2qZXLfyKUjYMhKQp1RQj9NSPhqRfPe3V1jnMLv8MNclM4/1yuE+HQWH
TNqST5kKVfeSWgVZJHiUJuy+YeMfjZoAVPFHZoh2N6vnV4/yAW3RgZAwnySffqOS
EfcDyKa7pFspRaoH9SlwYOsUXTBT3Mb+R4a9nkXm8OqjYvcXpBDMxBZjJT9ScSpo
pyRjmQwlJxISdwL2yDDwcd4eZvMOXdIA+RlRsFWCTHwgtkNFYYad2nvjtFnJI71E
xXRFjC9y4JI8Wh9hrbIBkhSiS99FpPoI4i4j9m2+luVXIYScQU8UNllD57n2LebS
lhZdxzLODyU3eXB1wvo7Z8xPhOfGdum7a92Vs9UAcfgWzN6rD78Ey/zQXirUnV2v
epzFA7o88DQQxP1LTZHem/Q8P7/zwX6A4mg9N/swAHJZjcbHstv1Mmai9YtLu9ZH
mb2/JthbX+6NKNY9yBJJ+82b94evluOzZD5YbHUx4kT7xjEWa5R4G1is7srmaPLh
jq2ZywCiDZs0vxKa5QOmQ0FkUgrm7db3903gflEWPS3BUDUsmWTU26QiLNe8kCah
3megBdjRgPHDgCUaRUfOAoRF0I2p7X2XxQNfpkQ8pfFbrHTklsdcTDSvqd4e/6il
3MXVfVnlMJlHKSmYp3TxW5uwGnTgYhlnmpURYmUK+iBh+oCGLf/YGpelgwxPDXJ4
YETVPMFEHy649p8zzAuTrVB5bhQtPtKfy4d217ES9nR1ZVE8ZkHrbMIGKmwDL0H8
Bhzr5YLkwqeVKItRVSxyH20paYooxDhGkMbWaAnJIHj0e21AnTV9vB4iRa9L2Krs
TVlm92+RUQULGOm7qkNaaqPjvKyedfANt5DkCD+HNypMklUp72MiUkXUDUWAKtQj
DGrvHjZ6+qQ1J5AUEsdQilBNL+gczV0lYS0AxCI6Als7jb+skRDDid57pw7CQMPK
LvBRPeaV8aS7lyjMO3scg9R/wDvdEAiElJbVNdL6qmz6oCBBynn53pojXCfSkZvQ
E/vGW6fVytsjGA2TX/pqr9t7ckonjZeEPgLNHQ0uqOeouUZV0jDpnIyyJXfvDvbn
OqialzvVeL/T2wHB/oX5mj1brFbQgZJmo1RYNhEQUiIOyn79ChF/CusyyNUumJvA
ZsNhVlzp4+ElpH23z1Q/WZPouDgDQUQTv4rMsIwFGdjgSCpM37L6xtkF9kmTZX2g
wxaIJOgoJbwOK5dSekOcowrOn0PNddrwnBgK0MHTSHjQRUwdavEPRjkSv1zK0we8
tRd3vWkzQJ+PgAoIpXHzq3K1SNCVEJRBBE50L08vDRg38O0Lgcvui3K2/HHajRua
vIvEV5grKTCR8X7zgE3b0brsdTWlxAV5JA0FAh+o95enmxbkYfdt3LhBYZQ0hBrb
Z/BYjCo0dFax/ccnD3mYqZ//FwXJ+8Ymufn201feO/m7UFz14lSkrkpFP/pBVgEx
Y0yrkHVHstpe0zeFO0lwUNS/5WyhvQj5GZD4a8pNhFCjRFh0LLOElIh1OYwyfZVz
IPObp5BktPgPV+Y4NT+Z8Aoy7z9+KVKWtexLwyf368rpmnE32DU6IxhRHPa5TjUO
vJMhtor/X1pjL0Cr7zPacNrclmU+U3xYkyvgAZBqoug2/SotO+tUIt3i+42FHeDG
iaMy+6+tZNZZcbLyM4mgNTdUzmTDrpPiBiwIyzk0P+aniib4EuKDfNChk8vKlUYL
sjN5t0e0gqCNkTmTh7tdqlCpWtkT2jBzfbOoiLjMSPnlaLbb1GFzovvbo17WSiQW
nfcBI2GYxhA2fRy1jBDVKtfxYsw+AEG8jXagQ4sMU1Cq2Jy+Zh985H99KdpSGj3g
VThJRer7Xa5njMjloFRLwCej6YeAE8YxP6IAffHQ9MilV1pp/ScxQpluvjiOP3Wu
1IDiPH+TQFdVBdHf3+eo/LEkHjZyOHNhcwBC856GYyjReVmDvysGRIIjXVvVlYOx
TQnHLOHPAjCRRdMFztzc8PWv/8FY3bU8XuBPOslnSjrUrDIxSu04vRtzEeJPaNs/
WD28ZokGBF4eomIAzHbAEQfUHHbi3r3px7PWgA17QKrBWENPy/wrR1j4WPS+JVcy
X69r+bVe+PCC7U3/81mumMqYnW83ePBlDXQKfyVoo1uY9E6ee5gS/pQKzt5srWSX
mxXR5AQk/QBjouW4omvgvBGFcogx60vtMN8w+3pIruSkvzbvdrGuCL4x9F3fRsSM
mK4RZDw/qMznY2WeyzioCZ5ubwRQZD5mPlUZD9fGqMet6khAAkqXqPhZfsQXSmuB
N1TTVjQgDyNgC9gQ+egow138kq2PqN0si7xVLjNkqr+V5BoN7kWVbK/1CRnwe0oR
bBvAAx9kkSm7NHIYon4fW9ajKu0fn/BeUo6mO7tXDDzdrsMnUH6dDtmkUrqrFqs5
GdNGHdYQ0natkn2Ks46lqp4AG46oQ3VlME4M0dKkq5PPUkmD4IeKdyYTTAV99nh6
gsAwVZ3BhcUfB0wMIf/7e7gWKfguTax54tYi888uR43UfegKyTnmRuqD9s73vYBj
dCDSACznNFvbL/3TAzXjrW0QvXfutOEdm6uLwkPTTZczvLVr0T5KJYx+MRYCwV2J
5eFXojbjHELr0KtiDtw5CpRXNdBpGzA3wfX56pf+fJVBKc3gp/XIC5j4O1k65TLb
j6m0qCWWZsFFOxM7PyKJKgiE4rj1JcXuCXancrJ4rxepun4NMbek7wegB0e+cpo/
1eFgtrn4uSB2ZGlKGGW2KGNauWTtb10kin8ok63r8JlSDIC97Fr7mz/3BEv/KkXz
q1zU32xfHMNiOGWLBdUEDykwfYkhGmJHpJmCRkOe7qsNPjGtM/zVmpWUN40AIgnP
d8Trpx/qqIV4G5ml7SSjq0axRG5/wsv3xMfv7Sv6FlriFMKCG65FG1T9HkmhATua
BybejOulHUV/JUwuswPtWp3ml2pEApPhJx2Kf80nepDWkEQzen5JJNbgqx2fCcFm
EtMailpdJ9UFtVRObRHOLTngx8iqh9LMDqVDiKgwpu6IbKybach34ZvC/rK6UUH9
tt9q9WwzyhsiiLQBhUhNHp85jw51mC46FQ/m/zzHgig2qOHuAEAsJ0T/w0TSSqoe
wG6zcQ5Rpz1pv5O70SZOPVnQ2+hK/+nBQ3Ku2eDRlBts9p00yVJLUq0pDaXoWqPh
wopspddkq0amewfL1FdYmsuXzUlbBaURTxvpB6fseLn4e1Bg9PBW6j4BL1PLPdRZ
pXoxvaMH8Qp7eYo69tEfeVMO7tBYHcHZgNmqAvBZW7BSJ2M8Ek5v8VndcQQ7ajYv
gN/gBxl6tePLS1LSdedA2i5HKbQwJmCfqtbgpTVaIAFo2EL47m/GHJ7KBiPFHH0Q
RXgTLTgj51pN4CcLoq8Ax7YajwXEDNzxhglC+ITpUxfBw+yxRkkGdq6U2BQ6XHve
K9wTtijezQ4hS+nkWDRwKs1kNJ+VayiKPSv8a3QaE1EWkXGZrHS1J6Uzjm11CQ0V
5xYPuRCJMlwkWrjEtFxVto6o3t9FEHL92kBljuOyeehR7/2OC7N+UtdieHYuXyOU
TpiO1843TpFlK7mBp+q5Vk09t5o5pBS46ANcwGb4du6Hx56+9Fs6DFYPLVRVeG9K
pkh1awS2yVssIP3is58bHobGXYSOhfmo6s8bdi5ENeGf1qHdZUh8dgcaovkj5wl5
CBtxW7FuL6QQAGQRj0npdqzE/JYNu4kuj6ZdA+UWYmx4cT/3YdkY5q7HsyydFPMR
OZc/h1L9N2jx61ceHU4jCQPArcc2g/BVypFn2Z4xrdtly8HISnU8DVvElnLzm2pN
rfg8Q1HHT5LG57SUwBpAkxXlt6AIHYtYica9rjHP2kn0Dt+lpBB+HQB+3hZm0uvy
5Sfu8u3zr573k7AHAjpYCzqI0EuX4h65RyyIyjHO/KrNi4NJOa2av5dq/OR+yYRG
Nyq+9zsk+CZ33wyk24BqvMfsFA5/Ji/tLFYSdQQxdYM7kRhycmI1uEE5ouLFGRO5
7gUQxyoqTa2sZXZhjVnrPlmngmwgNLl0wSTsE+gD9vF6v6pJ1F5yQa0tUo3+6qar
ORRvpIGvT7PIr/qwyMkPr700EegXaPqICXgzlWWTTE2kgmkLMc7pdCqYdi1tGwZL
hB/iHTnaNMhOty5kseCwKEAh7gtEp2JbCKw32m2OuPsnk4dWDSClk5Vt0S7aTI70
El0IkO98WvIBZIX9l8zaB5OtK+csxXS9F3i/95s7ro3u6L8T8kez6SPeDcHNuV6O
BBBIPG1bB3LekYJwjE5mUK3gwODKPgmEu02BF0SuC5/kp+SGoj1tzokhBz15e7xi
mps0flmS2Qb56ThPFr5rghie55NmTS94SBV8uLTCJvLVRZkwzbgC9I4+z6wzSqsJ
KYaja55//4emftNZP321mxfKxTVLetzWzs+bnl0w9BYe1w8oJsazQhIAlatd2o3r
TdXFMRuVX3+uLLBoHsefC63EXYfxkdSEnZo4HzsnfDKPKJ4TVygpDskrLzuSGLrd
Mvn35D/4eNXL9XSRlMusQkypLhQd1tUk6Lpb+M0++A0wDEkBcJ04tDDtd5VJqTZF
UnOSFSfOMfB45c7ExoH+ztCT2dFmVWSG/jlA+C0XI4OSqOvzFw99LNnd47+5Hcj3
ZZMdM4Nt9ZdTkS2ECl1DLPFQKDekJqFsr45/tws9GXo6n17dksjbxgH6hlX+Yl4F
1jfmalx3mhGNnvCyfVjcCeFq6g/Z8fxvLc5Z8bWwGF7fpR7t3BUva2Zq276cNXRL
tnv/qafUZB+Z3mzCa0KHPF9UBFFTX/Vsm9yAjgQHtry9pBY1VP58STvM2zDR2Ijj
Qh9r9Jug+mvY/NgFrTMlZIdu18ZX47GQSyR4k3+2PQA4dwTKU/4one6QMGA99W+i
UDjrJJDudGmlv5zs6KQWDN8QvPX5DJ1nD8qJZI35OT3CCOht4JXQR3eAMHdEis1J
78uu9MiELyO510HKx3xBsFOgt7bHbj6a1Wh8SirjWQF6ZhI9iF9ZK62OxNz8fn2x
OGXf8Om5WSFj5szzS/wO7PRSV6UL51U+F6seWoi6KlpwVsdLvG7HMY+Nni02wPqr
7eecL7Vml8mJ7hETqpTUAVEXbHgXUjSBgw7Z/I1lXWu5w7Tds9yUhBrCU8GaQBRJ
Cu3l/zN9SbuKPWNC5ZA9+vaRyjGUZXk/1JAyZjXuzO7UuE8IivdgJmirOIiy1edW
WdWtdf3sATugRTs16hgMsKx1Rm/SCRiBvRaFl3NizGJyfXZoRl2buHRS7lzWqLd2
AeqMPlCMedQY9ao2rsSWoxoWGI37ZQf4j66SxjWQ561n6/fh3/o6wUiaFh+Q5z6u
NFqlvwgl8AeKs5o3EdZR9uGKHwz+29EZVnHMF5eQUmqg8izFvWFq5BuplPTpJmdR
3dZSpIXrRKbHz6EnYw7y2uA5hSHVEmUVD6/tMWujS4kiaKHZ5oM+3UvuygxzrZTv
m4dbCDgt89FfuBt77TI1jCKLrCK8NQbO2dPltDcWM3/xaabaFKLVa7c/uHk5BP6v
ZFTcXIFkQDigtCRXWBu6yK/7jTiBh6dVj4KNWcF6T4Nrr+snaErsS6mmkm04+Cg6
5jpZ4dE+6ftcd34CRl2UYbts9UUzapBcwH3JkZR8VwybGdu6DScnv8v7yvDptBYB
Op6/oEs/KFkvD/4CM3e5UEqIg/rl63NVsiAu1u+ile/Ic4qFxhM2fwPL8caHSxG4
31KBFb0LKeC8O+M2PvFe4WSs8YcKnj/sXbII6RsWQM8r5kVipMnq2e+5leS3C40p
1po1b1DHlQpMPQ8/HAMEnicNzPS+6IAZ5eUSgpbGER5yNdcmT9lvNQVvCByZsPoh
46RmADnpLxr6MvAtHYvqWDXODHjgtRbMqbr3hV3hYEqJ9NA3U3NSR6wSkKKWRyGk
1cfwlncS1I42SdVJmND07nektCxWmy7eOH92hgbx599Ox05OzDyWlwYH616/U3T6
q6gxKYQc65hhUwMKIQgdsxVd0EihjksjT2K+ULjXqYDsNikK/qB9zSmm03m30m9J
1mgNujYG2FvFmiqZC8lQOlmj5JhVod0ly8jjmnAz++XjMj3BFTVDCYAEQ/wnqXbT
lhFg4zDl3WI7lwJhM6nhuoK74ZVzU7EwTI1K4ue+LzE+jtX0bXSxkARiW0ZHYEJU
dhqV7bYVMybhKyUof/QN0NFXozdBJtNtRrhYwWmff7d7QDaFo/JOmzk7aVGkOBXe
X7ge9K4pt1nz+4UrVIHMxXCX3UOrXS60sIrYcLOTv8bXuWABPhvx+Hv8xLuwqXHi
qLMQTJ8inrsnK+6RqgZQjN1Hx47OJH29qj3TkGTYpVrsPwyzmUnkCPE6UMsHvIgm
TrrTNPAjEcbNddx6UTzBbaZpCvPRsg+26Cp80dPi2gjkGV7J4ljqh0lSMefjiTUp
KunyEsJcpBa+zZ2i4w1dlDOMM6E87+3mdKh8fzgY3sB71dI0BGzFGTx/lf2p7UNF
FUVTUvUBEu0MjkLU2seXjdTW6IffVPOP3H85K78iWigpMCIcS2UH+Vm/37lGK+LT
GxANfItRIuAAYN+SXpU45ahhRtsi9Fgzgc6sbt4Fh4+Ont/oJRrEzDNDiNBMvNTu
UAT+ZVGi2bne/ipouSzKDvmyRhnSONEeRCT3WbklaYM1H/SFgGF6/bGAgfSJ1ESM
rfN/uSeH4lQaJYuddppxo/Dx/ZXoQmsgnnukGLV0X21yJPqh0MUkP7oOsmce1p3W
9qTbFllrgAnmGeOBE1Rk3DxOZ8N8Q+Tn1ooYQm8qrcDygZ+9bwAKTPxZpqtGQd5u
GqKnVCr899ABAERxK5pXLfykeNaeo5bgQYg/sPwtJ6TWgO4LEcH3/6PPGaDpkNQB
UCaZAi3dGXB4OqmNSebWabmFN9livB9jYMEqZXGiAGIpfI9rcut8bcE7MQH0XIxl
fk+Pft5oCZU5PvGAztqrTC5Km+5JzXf5jHL8WFtdhjpn0/nTr6hA3n/ynAldumel
S5qEl363gWbGV8rziVsDdcgXPjirO+nWpxY0rUAP3mRAMwskWZUl6t7KupjTQnE1
HgldWvxNcRp7GgkMUmTvsX4kc5WW+TMD6fMNKNzG0ADzT2qYKx8hZ3ChB3zyU47/
IjNdExbXR3wOeDqglrwSSDh1ea808G4ApdV03ty7BUFCnGXpzgpUOo2Se7UPYWt6
OeCyisnWW3EKrpCBnK2lqrR6maSbbS8U1m875VVNJKSQQyA5Oy1uNw/n/s5eh6vi
RlAuaXnrMLk//ZU2w5tBOh7BhPJdeoLRzqfGCA1xJOubETQqMkrLAKpu0k8r7+lb
EUF98/tadjWSgEXl2O5BR8QPJdQnk2rJvqn2V+zqHTYYxwgm+49jqYBet8yNskOf
9GOwn5IfTFY8HglYNUtZMiW1B9DJwCPPN1zbQ9CjA4LRg6AYSrlplBN9ouMAryoq
rW8T9zOPAR3YA/lvTKTwmNGVXmYmu9J4MVAgoiZbANCjYY2Lv+Jxd7xiL/PtXdJ3
/Af4vCIttUM3+nPohVns1hlUhIGGOqXrfa2+SEHxW3ArXeCLVUQPyyMuObhIFC8m
28LtFcI/M8x/HhcAbO+Y7rRvRJa6XFRXMybr/MpucHUXGyjK0ntFJmlqRqG4BCRV
EnM59lccp0Uj6UIdT1bV8A9+wCrMbLkO0mBWSF5qwrBK1g93DSWoQa0GYBbShSf8
oX1LWlz+zRozy1JLIIRsCQ1x6+ts+8Ss54og7tQkG/cwfuJ9wf5+TIBA517pg6n4
OUV4d+MycqRvCL6ln4KrdrJsWLRoMEz+lj4cVJNW3YjIdgEq/HfC8S3sOvXV1FwJ
MPGGKY24J1e9DGoKYgLNqtAv0GN7GInQsGPWjy6khqBzlZWgSDya4/2vjn35s8pz
FlLL5nxgNhByqt71VzJpaO0uCo7wgoGF4umICgQ3OCSKo3RnYg9J5qWq5SyCGh4p
frWilViVY7RXno9UEFIBviMvtfxyIADm6KB1M8XX59T5eNpVk0I2l9CNFObqVoQy
oUUPPfQ8jjhDrlJ4oNtgzstkqwR8Mvn0nkGAa7g0etDQaTYCGmR9iDwXhdFV5Q4T
pSk+i5jEihpbbu7FDSRfSW2PxmaPdRvpPFTuCSRZMMO6/B8h6ArgP/E0ia9rfW0E
RTlMVaYvpLhIQpk7pqqvqxvLj/JaK/BCtjC33FtTObrm8gtOFdKqfiieHIJ+5OdT
OES0A49pADS4kXFNOjZHlAlKCo5yH5z77fEYBnJTQ6Cf0uptX7UHBI4bOg2JBIbi
Isj4BCCoHBe+p5/ZHrvAI84aKgk5jJsvHwAe8dq1vWnCmEmfxMG4ouyAUyPCKBvE
CcgpHs992edfDqBubddXJEYbrCIg7Ivlu4qw54dnoNogSGTrh3cmkgzWS2NroPEa
XBM5tW90/n6vNv0qj3xQ+LqWGf55Dsw/5xzr0ex11AjvRtWxMrPyVq8FV9p5nnsO
/VRulLntdnQK4A9qTd75ro0p0EWxBr76MnNZf7ymm7qnMsz0rsQjLxhtvXVug7fa
RMwk0+65CltZqIu6G2bsu/FHyWCh2gALtAZXWe2K70Y9KXkyzEinCu5QsPIGPBWD
7RKf4s7hK0V+/QlA+SACxdUvfQ+nPrfa7b7tryWtI0G3lLkthnC5AbVO9G+Uh8gX
JyQnX5zHAiOIUQBspBm7SlsFCYt2nNglHhpswvH7fWSgL/MqxlIjhzo1vijw0/tV
KylXGgydevMgURJho6jwwAzF/bBaRbGNQSA4jPauL6wb2bgGAF1tklC3aFCE7zxz
NEA5k+HWF4OPhxt+kBk+s83dOcDaaZbkPE/3nES49ASOM9uE7euQ+0OpWaXMbCTk
9ncq180d6h9cjzg94f7nIjtEOsooKOCDi3wKGaBytx5aIpahj3kigGDc4Wlc8GIN
kNswpPcTjQjSbZYHI5DgwNXbtMIp95/EbgRnR6hfP1vEOqJzZj/H8uQxPPbvX9vl
LvUnpxWNHYhS93ww0z95sYY3ErzUW/2qv2FKtmUJo4Nfu4ceprMway2D0Vilv0ax
koaZUXkU/Uc9IAqiJHkZvZZsqhQO5sTf2qUQ0PhXwS4+dtwQQGQwOoT/OOs8vSwG
edjru9zbzenStDHOFtEnhTUkxwrToaVSMx68lU3dHYbdW2n2wdEDAEhizReJRzOx
h4ZnYAtb1Z0cy2hP9ssS3+4p8cmDIg3tZ+qijFY7AzIxD8F2ZenjKL2XQrfJiNKc
TcPJ6p6A5EWBeIvikFu5wiejsXwfb2Q+wWUlsyt7BxtK+zQFUT74oFBgejsLEyuE
QJVVvhgJze4enn8cjYSxdn9aKefHxwu7fOGKgydw+Ek6VnrLwogO4CUczZq2i5OS
JckzBGIrkrH3cf+lu5Z3GAvQo5kSg+emx2QP/7pC1jeWfZuS+bZIvEO81Y/hqtgV
aeoXpVKhW4Ryy+cLXX5N5Xo5aEjGNMvkl33LhiJEXOr0U1l/t7R3oSMWRUpniHNm
OqfRTYIveIbYwnMTY6lGaHckeWe0knie6kiKQsxKykGGpCqdzqWHatPVcoBMXF5q
HAiQJwRCkmWiu7C7CHe8Y5qedGdUSV+u5MhLQ8lpg74uEqoNrGTgcfdtTwlNKhsY
lA26aMA1OnWOcH6Lde/bWK1hqa2OgDQZbRVWmNntIbkroC4JoEKwnwNrMXmZnJuP
sB2H5fIikdct2XWVBbUZngyMUCCQ1R4R5L9wxy/MdBgixnR1k9FOmdZi6w8S6tmo
b833qmS+UjolKpfvrkZQjFVrLed3v3mhWELfSsVODS2FejxRIEOV3y55SycYFE0h
CJokG2D9ACsQ1SORUTFfKZpkzb+tCx3w5+HoHv2G37bfCvSTxDxQiNVH5pLm6bom
wAm96SSgdjh9sArXPLJSM5oU1xs1eBIrfZDQtezRmM9qDOwzIu1xQrJz0uls37bW
D3cap15dqvHTOe+AFMaRzhaNir4UKSnhLiDoIDK1tYo617dcasqzTuHyJZEdY5oJ
TWrO+SmBm37qH2ugWGof5OmyNqbg/GRJYTY7u6sy0FyPsSW4NgPDKsbGi3XfTq7e
uS/KNOsVaw/5OVsoo16cDs1x37eeDeQSdioQ1S/tNbe/1Ivmxsc5xDESghA4loK8
XAj9OCcw+Vj/ERcCmr4ugLR9qvib5pWWxATVScB4K3IZHFq2iYuuForAGFnzj4ea
owyf9A3NgQYgZDEsYg51VBxMsLwEzYABiESkz4nHEzSHaRX4eBgj5pi5aQEyvzP5
hKCZctKItogx34VGwRbsobD7rpXl4JprcMTY8v93TA3TXc/l6t383Amuezd6O5qi
gA8L++qtabLz+OiUHRwe5/E5JHOSKXd1Hak+F2yP9fQPNPZkHDBZDF4fFxVOOQ7H
QjzsxhEmdakvOfQZHeId41JVB3qfcWpSNIqjJpBOewE9T4AMaY/pCcmuSonZ2ZTE
jg8NJdS67x+p3gRcmXwGajuYy2piBxiGIjFNjVI0CK5KRUusbtIKhTz7HF+TYVUz
8R4CVrvR3Xu/B0PGiXP1QX3K856hIkg/xSYkovy6guRxPNcfzSz56yP2G9EnHr0u
lJCTTdn6tUCTp1aPpWAPR/tfp/FxZDqfu5F/ZLlXvieuUBMvr/d27DSTezkUddBl
p2uG4G0KEMd+xmwBAnFUURfzMsfuuOxbm1nbXQVIsLWuEnyTf27sVMBzmKtd2qn/
OlesgmgnBeawX8IEJBdNs0ir0iJkonE9rHD5fEv5kiJmEkmuNBBkZWftJYkBHFKS
eEwzmV0G7NBe6uQcthuudhqkRmO0YD6jyfUez6VuO+5E7CPNbRGAwIQiYytqL0vl
E52s1PZjiht9xwhUmp8DB3+w/4/d9floY9hjFhvhFLGknVPApWrlbSWEIihls5HP
NQ8243NsaaoC/lglyKSP1CTY9sG/UgDl+/QVw3XuaTOBBJFSg6w1ehHhEqRVrdDD
J+bg4doa/3NgKbnadreARPaEyoTFw0aZ7/7RTMcuObcectG++OwYiSWYDGsyN2n1
+hyEHzJme6EsamwAzcJWeXiYHVNbN9ZFVwlfK2DFvznbVlTpX5KWI5axnn7e2xAn
Nhmv0DyS8BdD7sfyrqMKkLgqrvTGzOHGC1kU8ZCYJ8yrUT0ELL22j+d+fXaLW7MR
EsB2FQV9wewtspKX9kY2W0ouuQ84DSKywc5Zy4WP41kEsfsGMwlrh+fNLLxV0iiC
9rwESowVpGSfdw7Ojx6l1UswBCcCnNtXkLSi6+OHM0AF7KgBlQ5zAh72vZCMWENP
ZVDvikyRA6NrOoKuiMxvK2WNnF66Jse5pABtkddwM8+seYZ8p+pbB9AHuOJOYZ5D
hsCmznyo06KOCbJwk8fTiVXYTpHbHM8/Ef2w4O39OeMkm8oSH/mJVipY+tPhF4My
cjzpNimxv6ngf14EVCG9q3hJc66WFq1rXggPYOy8AIXR+nsyTIuWu2P45mtq0Hwf
Gll9OsZBO3qJY08edqdQa4Zpm7b9Y4IxhIxAUKGyyX6Fyz7ra0jY56Jb9Fbt1Jp2
x2U4lBL9+3cf3JYBZO3AdPSBZpVoc3IFX5updjZ5ZcBynblxB5BZ6lnZbl7LMMoC
Klv1Q5XEy1xaFjQzgnsWzXMvVP3v/fSFT4OGOhMSj78dp1vkvAELBKtI7yDdhFYm
+Cmdegmlo67F/6MkRVLOALLE9E0cu67j1ZioNetQHAruTt5vY2nv2WkMV+b2UD56
h4xoiXdOiCEjgEpz3wptFt2VCN1wxViGyBNnmMSPgfIXFecmaCVOkVKAVgl7Mpzx
QmNairxicqWF/J2zKIPwO/i+LlmHSoCxz8Gbiyk7ZxYS0Z+QgjpSomz9DgeJSZRS
pc4nF0orBkEXT18kQIkDz1MSk+ENsG+5yIign4y4rpM1KX1oxRPa2Zl0EIMTSKLm
+beyY9ubl/Uiu36yDfbwJjtlFPNQdyGKww55SGWoWB7zQji363CYXZMN/kqLl5TN
urLowuMLJWIbNisjI4b7gopDnrFw5JGx5e25/M5vkFlUeweW1xKSRwFcjbnLP8gP
f+0h6OPDw5aTeodytWX9wlvzruA3z0O7qYm/pFf+5Yd5MTZj2cq+d9MIjS15UlIa
TOlz8yYBxtESlSQ/NBGag8tT99gCXSnjPISlkhF1cFlVcUU/SDsPS26jg1u1IdHy
aA/LfVhi80MYmZNV/A/xiMKO6ZtBnJIKR0CXZxKqNkHpKM0EeP5CysgOvy2h/fzx
LZatn7q0ojQPFZJn/XVJMIt3VmLyv7QizDlIzGTa+0sRX9KyKa3HqUXjOkLn4PfD
LmkAD7EhUH/O7QHR0I/f/PXv0WNLCEbq+9qCqPbXv4VINiYkqK/jKEhOQLCPQ679
rIQcO5/bbKVicRTAFkqRnTBp6DDsilwiYouOnn1G3OFpnHED5TFtZXvQOcun7ncQ
g6MaBSn1zU1H7SJ6VZ3wQ7isKdxS9d4juRoeE2QVuDRbyNuU18r9UuMrHZjPCSNs
NouWsLVX4vP33ysn/IY/lw/XTlI1VuDOcIdEkeGaPLMcrkQK4l4jrnWF5Ji5vwi7
5WXMocK37pqTTNqcTov3Cksp1mSDElwtFuIhrYk7FiJfyyMBrYrriE6Kd4eCmGpn
Q6Zn2zeZ2pbflka+bEpI+xyONee+gGr7qO01v+EQQVUp5gdpWCVfabJ1J4inFjL/
Q91lYp+F7aDyVC9OLM4cRLImU6Nf/e7XNpn5cPmDdXONp83kdQP+CxLTY4zKd7eo
oI5nMp47Gd0PI4U2DxissAkg2Zkk8yVn1sjtLnnOTET4yigMX2HD+Prwg5uDUCPF
3Tb/EjgZeNvEc0b1aNPj07Nk9JGIuV1+S6UqDVqyVoV1aKtTb1hG4uZMy03nS+kK
dR/x/upUjSvb0eP/s3NokXKBv28wZOQz48TKuiLllBbCibsa51sQwpUi/xogW0aw
/Pq9P2/lXTHE7k8qSIkDYdJt1GFV/wzMBLYHZzOSGzFqdu7REk6wqE44qvMzxu2L
wsoqXqSV18WSXK2l44kRJH0Xzf1TXrMrJ0BLjqYo31PDVtcYlcZhf/TImZ1kolNg
tpdzwUfn14BfOIgt1ZIvuXvp8xQ1N1/vgewYL2M3eFerRvaEN/aJ8xu+AG6N0qTc
mBTRznK3Ck6HUHkG+t1mECVKruar/Yd7yKeT+uM5F9fPxQi7bUY+M/Xnlril7LJj
1J8ctyrmYOsw7V12u5wOafHINeEq2sxVuQoXqR0/n3dugjGX7BQ8wHVsGk+Vd67X
rMRY90M7Gh2TEoNjnEFeNFV31DuTWI3bQmmbM0K/4DePNN2VvIDv8I5AcPrBqMlP
TSvqE+QAeTSNTegpYzH6Z/KkHyj0xVM1LU+6zFyCemLwpjFHsd5OUibGOSrjyGbt
P6j/Pi7ReesTdCjy1cQh3jVwy+SQ2GXTSEhdtLr4SjoJhfpops/4MLFOpBgiylzu
oPGjFMUEBgq6p07XSXug5id8jeDNGsS86LQwY0G/M/OBt3CiVscPVUD8wnx4W/yn
KAVJajMfCNbyev59XZb9jEX/wWY4MlzXxiclteuz9Z8pylIewDL9XNgP/2w5zDLA
4uz1BcSlv9lKvm/Sb6OyUBFHMQzgoYWy0Ht6v0QryNvsTQRt8Qk9D3ypohWvPpp+
2VM++X076Jby8juiKfW9Y+hnerI4CAQIGu/jUXak/a1PDecDvB9fDWmmBH5MBAdV
wymHg5iGfavwbDOrFHvsdbfYudf/Vp03pgFsjdkk+ZaatVjtCPfLwsNPPdqeV+7u
oQokM7XBxGxm9x70HItF2AAYDqXGIqxF91+1I85ybwrkA20/eVwarZEinwTT9VCZ
Zpf68ekTrkBystp/84WLl3kFRsDM7zHdQUoCg7BULyFjpaEOg+S7uA7wRGih/Uss
NOo5pkhIXHhTmXzVVyIzJcKGYh+FHtmCB8zEGklKavkij919wzwQflqvk1lFG4zs
/xILBiFxzHTr+7Sy12MmsAS/s/CgR4oNhU/4n1kh2On8aHsmgNyt7vLZt+dZXUoE
UI9HR7DMvbTbMPlOVxk5MjOulrRcFkq6Ok8E6LcHzAR3+tecMda+o5Qgg2HBkiCu
Dgx85hUcajBz1LV+HGEtbDlitWejC54E6WOasiQ3A/Odqt7yac8XsdPITflkaA/m
Mf/cGyxMsgSJ4ljWO+zF8uYY/WgcywyLte+QX8AJsOpit1TxiNxAoPj0SRGjzTUm
obJFPf0Mc1/dat8oP1APzYVyTNwxAJDDPqVDAT5HplthE6fnEtYNLbnHguW694Xt
7mfGGfYLpHvjNIakNJnnIKFiFWkvxKaLEaZAXOemu5BudiLrD5BOnTL2zHYwB3pt
8r9VamNkFJCsK6S7VJZBLi2CJZ3QuTVXTC6z5oDlSL7igukwgdilf+9Z8IcquTnC
ofrISak1IHHlsmbatkiTr8R7JxZU5lpEbBaAgohqicxwCoi7lyRppGhO6bXL3NN5
j5AdPc0mWlcglHjBz8YqJNEuAom+W64M77upbHUhS1hIWf8Yl1kD6FN9n6Kmpf27
0G/NS51Ot+aYPOB+4MjNIcvlB8+QanxTBsvRLx5h7Z6bSt4sJHT5LsDqLCyUOW0P
hDZLAljJxTPD1PlcBsIxzrQRXT1DyNxiHF5FSNR/c60lMVHo0uKsQD8RrBf1etv/
jTo7b+yhWwe72DppsStp2ZJ0Wl9NJpo61e9YKTAQhGoAK7f3GmkG+O8DTOKHhy7r
AVpwOvSZUyd+O23DKQnuJidzktC5h0v9BqafDzFztq6G4AOIGi4/s6K5+Dm2KvMe
EomtlnS15dhGHeYFJicZ2nYo5c37RkzjSg0JpxNAMr2+O1ZIBXMOBdUYLaqvDYFj
YwKAj8YdNbcGrybll7bSjGphkd0XKka/G/FIONXs2OMDJ/qucGMJfGTDElZCj6Qe
JeW1P+GbCExT0zi57Mj9TxmedE3JXhbs4FxK9g+MbIbilDP+2WpwoMKX1x6tcdmU
7p8BaWvjxehx9+Ho7HRpoGt18Q2aF8vkv2GViG4Q5NuUgqt7T278fE27Q3jZtDbt
q8G0LNY/khSNIdpHkci7tea1TCYSgb8EghhK/ILCMvBJG2c1eewarB1TRGAiBXTZ
EJSdpwC+73i3BlrX1+UeNVjy3za++hdS5C9gwEK8tKA8kML3it5TntI94K9jt4s8
s+4GyrJCqu8+L/oYHuoZ0bax3sdCfTPC9XyOJcxoDZw6d/P8iRam5StKSSg1CEEA
2iCGjgAGiEx2L0X7dWwtDIM9jap/j5+lTIIZ5zsLVPt/66rKDxAKzbcynhxwrP8b
y+LyZhqhiiEcI/11bfzIQgtquoDfdC2+U1Hg3ILY9EMvBG76OQepQdA81NdaPc3u
daJwYAj2GCC8Uy+QyD3RnJawnCcYgQ2z4isKmQSf3yeYn0YSFGn3/UeHjDLHWRPi
IWlTpDtjBTG0tV46J/L6KiyKtfpXEsf3F1151B3SMek7q8r4iZe73k8q9P7k5rNN
KaSm2JluKzY+0GSKusTpoUYvTtaqPUMUL0Wo9IRUfsF3LFScBu1qcrn/KFymSGcG
LQpDpQSoaVWmSmMApFN96kF5dXQAuqnBtnggqKuV4QhIg9uA61iNtHbKv33z7FOs
Yoyo8aagoyAVhftCfn7luhEgsCTPeY83LNpOVCsZX/awaWSytr4l7DDdkofVtAMR
Hp3q1yxpB2Fi933nv6abb+hqWkXvJULjkWA6HVXXehvoRykS+9qz0sRVwhHjFCHC
ChktJaUs1GRppLR0sIpxmNozN7i4eQQNDnUbjWmRMMc51pSlZ6gQhvykUmSzY1oh
wtEAekN/bsytKZgdih6MXKo/17g+dpQhtLaPwtayDGvKsC4hPXnfcUMsPidF+oEg
2WCdp7cA4WzN4zx41Aj1OSdPtMAu/+fJBUUtQQOwdqkKXLBHQWjVxyxpjusi0jIE
JCfaGj+JaFL1kIT+RJdEHF/e80s+dmBDrCWT6MwTsc9rwU9aDIrYMt45SkmAF6Dp
fxyHb9hDi1XVWQQJk3gStFKSI8LxRdMu0oysydLvR5olFur5DLPDxhLq5WgXF2m4
Ll78U/Pf2/7n8MV7BOfm6oTB0qPt/mgeSKaF8sMSCo81ehvcEYsgdJuwdWY8uOXR
OlPd/H9DLa7qnZEJwqC/cSgTsJmzY/SFLydWAzF4+e6DwEA+Cj+U5w5osINcs8YA
Ai8ZRoHur1qGH92mXVAkMEpGczLI+YYHuT3QRh+0OGf/7rMQjExYlUkBT4OsLWsu
uvMFRna/nfeLvbXEO3JwhukEL4C+WFxL2IYMsq1FmXmO6YIB8yYPP45zz++nivtq
pSlLJVJH051lLIyJwRVMnSAng85ahoPNBrSM26soA98XXqGY2HhosPKQtmO2NUEP
WexYMQq6KvbQmWrsosRtJWu0iXqET6s8C4m35lbcZ8XYc0NzwtpJFnY1Hyh0O1A8
mt5XRoAYJXFIz/89d7VL+Mf9HxjdeboYYcERabAm5MjdWDrNbIE1vc8uM5weWlM2
BEeqMvGEv91Oi+UT6Mx/H9B83J7Y1IxH8EBi6kUEAAwPs/epHUguj2vv05wAP3g7
iNavUtnDWtWdcfr7QZLbHXGzJL4YZjjCDXFOZ/a+uh+KKDmwsx6g+5BHSWR0/D3z
1t4jLJwDfScGPL7zIbyjxtgr91wHaL2cUlbl/uKn1qWFWEXzXDqBKLvFd9k5/PlP
1Tz/Tuh6W+Qrs+A4nksI8n9iEjINDB7ZLT5mz66B4ReEetH8mclSW3GJA7P/sl17
txBtw+7rAcPaVhEOFDQAleLZcoLAmNrqrRq5A7uJ+yxWI/TiR0ROFFfry2tvZA8L
zOZBzpKT92l5W4tFTsAjbrhQpPGPYq24RYJ20q56LINa5M9B+HvWfvChmtW+GJ4c
2vKH0F2VC8C5dmRn/oZLWJsJ1FuOrejMBdobDK+p4M4Gh5dV49WvQp9z0E0AetY6
QOskugSQO/aIsm///l9uNx67PG5DR5yXeAtQlQ7rCxbkTyT4BCnbpriaTbD4lkkX
kmGHIWFwM0x0bVcU79csuWP0FhP809JovrP6TBZlv97vrUNGZEDc+3EZSMgnnVhH
ReIc0WBRB8KDEvyORhkgTgpkLuC8zmz4ne7dfrEN105J+BTrW2UL7ZYYWtfPRHAk
Oh4hx17/m7A/aD8qdGBVWunsqkvqc9qnJh7gv6cJGfaNPNVBDS4jgZJcPOUDS9aF
/o4V+JSLx+gp4dJxBUvGNcsNz6fVIDzvohmzahz6Y9Mm5w2n1ea6m8RL6HOFepSN
bmtpgAcO6+2IjCi8zkO8JJ8XyIBLklEaRWhhLl2U9LMY+6JPYDCUciBgEuyRw/gw
hIMDkC9zojMnSYAqvrrr/ilZTKuqiu6H7X5KTYX01O38kZkSJmUF8vgaD+5rp8Er
HprFkedEFGLDqlT8k/6tZESlt6XiXfwHY89CXUhX2Gd2w6p4eQTlyjrAD+Q9U+7Z
5y4OtF8wWFofBHc84pHaOKil8GAoNQ4UCPiqbwixYncY48FwM+oV+rguH0bPleYT
pDam0VvZMXPvvPV35BkBJxHowWS3PNXEZh6RI36UF+yiVQUDj7H2NZaL0gbLNHgG
ZJ7Cxr/1pZHRctRp5oo5nK8a9ppKJz9+b7QnuYfGhgxcaDumf4qFs3wkDYk0RATH
2tdKkUfmqgZ8PGfmvWO21HzwP6yOTbh2xSOx9iryw9LF8z0n05X2IOGhN9xZYqo/
QbJZQNo2kLirpaoDfjB8GXNx+drBQeEhI7u/jO2AH3DaB16bxwfH51QXPRcRSOtZ
8LN/bRbfJHq6PaPX+JSsUQ1E5lDHusGwvEGaPep6OvLi3+oG54emWfjpjQGJSg7D
PkBzCIeUF//SkPOfZrDoL2k8TGzn1+eery8QiFeIVupIqRCRst1pXXt3I3JpnzK+
x1Qh0zizbRtWO0Wr63En9wnH5H4bIIQBqnOSx6SwQsXP7uP2zq2kRJSGmB24DeoI
lssQF/rDfz7bOxpPax/t6uZOn3ujQ/3yZZzQy5hf2Zq5Fx0WB2a5SqASnb1EKVcG
8zdMcLAVqlrE9u+83NKKgySfFCQKtbgWJgCdaxd5rrWDMJLUpHZt3tosYeOWJQbx
xsuJAXpTE2UrO1osqfS/diux3pqKDRykAjGRgb7Ky/MjlkZ2MNh+cq2e1ikG+qQp
W5ix26xz9Lg36m9d+F/BHlxgY8Mrsxd3zZiHT2xd2Uu1Lmq/rhGay07GVTB6u9qp
J1BVTtxh87xUM2WL0+/J9BCYz6pbpQvAPyGw6e3I6fLbkrDs/0rX1stq4TvTPDUV
pI1kVVoLJeJS0poftoHG6m2iA3uYUssB5VWuh+h0waO24vLzwPMf7Y9CUZzf+Jy5
rEY/dXADto9P0oWDuqS74qS2ASjfrGPpHFWR68OfhEZyvXyHcBiQGdJV2eLHjwkS
tLpHgvUM+K9vWkmtFlGsx0NJHJk5JOwRTDHX45DKzpXWfBzHJVebiAcC5SANM9Z+
9/sxxMYTJR2Sukse62I6GVXzNe4POROJc0FGlvEnqUCP53NVmvp/7dtgGvKvETp/
AFFvnOqgWG2/3+sdJWfG7lFMkmgYNOSNHMt4ESg7oO5XmRyBbZ1RiS0OPGTyoipQ
DFyZl8jEHL8jJI5f2TdA2uVfSgPYyl6mrZ5O6+f6biTZUHw4hNM85LADy3W/n3tD
LcfKq9BpAy9zehfaPCNvU6jSlQCwSCqz/VZ3MDdY2zv9ASRplpvvpGDz57kFZs2N
r2XlVooFEwWW1a2WVdX8G7Aoodhp34B3K12tyXhTkAjasLuVQoM7X8aHgV3X757B
YEmrXbdL4ZAtl2cI0s2oPv2pg6TovowhWM3dg5rP4K5YXzwmIrC/sBJq39GzrbfJ
FzPdn3lWdt1sgLEE+HD/VlYKSj/RHgVfurkHjDzbSe5lppfUBMwEYuCCJ5F42fOV
48oooFKS5g/WdvZ9NR5i3xFTEUubRpJtPO3ChsT+RLRMTPaq5Iow6e0OEI9WdxFu
F82woG8r+Z0g+sIkYp81+7CmsaIEjapAuxROUKEKje8338xEtVaXtaIlmlQ4pM2X
C3FHO9X6DjSYpjOMOfla0cexJG2WjmMAGTDZdVXUFq0rxTtoU2GirH/LiYEh/Kx3
tGviZPCs4UsS+AN2ylDb70Wj49zFtS718HE8BUZKcZEgt79bOos7+djtV7WnpDxz
376iC3l7kSBXNQFlkJBmapmmewvAVpNFXyY65NgQ0eus7tEFcB4tnMQb8QooVXZp
w7S3YZ9qSLcXV0n4hcbxu+2PEKtC539b1nLT1xwniKPrHQDQytUKEaanIL4uGpH8
PhSdq+Y/wZhGaMxP87k3ggc2EmJXRFka2KjXEbYg1p7AUfgSGa0tkDTzcpnW/DXH
TM65qfHxJ53lrgTKFyEwdT9CR07aaTVlu6vVcPaTtJlXCUE1FQXhtTP8gU32YsB2
NLK1PPq1Fe3m/btifoWYEKo5nrwwWo46vpX+uc++ynwhYXJEHVsmIY9D5vfJrLB4
sJMOg++Dw1kGFSNYJrt+6ijiFSRY5sHlK4W1CejMAa3/p6WGgEdo02EYGWwiRk4R
yZoTRhLwbCrQmj3HMMleIjnB1DtyFWzRyQd3r7LIgqAW4f2fEwm4dSYv/PV/Aw+I
SfIsRDsbZJ56nTzkvz7Di6pT+EsUVHbkAPPMK4NcigvHhmFEuMkRXV5nogH4d6bE
o353mB+/+/mP4BusdL2HJDxC15+X0tzNzfvoaZdN55F1Te2RFmMm/510LT/bqsbX
ydjFU8yrpuzOPL+f7fPj064A+w7WsuZ7zVtd9DXsXwpB/ALGRsAYsvdNJJZeOlND
QCQ0Q5knCR6vkkuvn5vGII0wV+OdmjEB1f7JGqXX1BCwO2hKCeEkPpYc+5WmfoU6
gcJCm+UMXecuzeiiOj3nl2G4ElRBmZicTLuGHVDDZKGrsfyAlQGxSNtU7miReSI7
3K6/c9MAs9diqFayXYn7Z0Xaek5PW101TTUWlzsOOFNIyxmYCIWc2ICoBG2bVqp1
io8NPJOBJXT8xNdn2CMy7MPEQcL7T8KTiwa5JGhbXi0haDKvC2K77NkX9HKpt3QH
JyDYT8PD3Y77h+gxYIvryULt04v1+W6OiCAc58CSYIEeAFX0WJVCJKri4NtxxyuZ
9FpaFxuiVHVZR03lZyCpOAUBWeees/fhz2LEffpXoGFyF+gTlL1/QD7wxGPsFbPb
O8Bf5QbLs6I+Db5JwvS/W6QVFEK7INPLo5LpEn1zxR2GufR3rAS4hPMdIedCoR4N
hwUSqzHFPlaCJTa6RyqsAI3eGEkhOkyJdr9ezzf6x+IaIWj/R5Q0OCqgq4cDWhzG
uy3xnXpwPYz4+LWmg81reJS4QoWgXOR3c6q+m/g5moa/kJd7YJb0PgbbSFZQyN4l
DiGjwUoUnugHI7Hcj+vXeSp06WDpG6bb9UNMt3Rw2XHGxv6F8jXRe4ky/7vBbcz2
yz1weWKsgQM0kj4siIsQAmWL4q1TnT3097uHZe5OgUyuVJDY70T6RThTvq+vQfEY
yMUGNOUu4LmPO6xdP2FGT/ez4IvRqFpc4DcGEH7ZzmXYjDMmbMLaKCdAl45AvWhY
EXhujRZ9gBFamrCqkLqM6XrubHDs5nx+62RFnMvfgYTWBTkkqu9sNJhBfAR69J1R
l9WMJOsNMzN4LBnzLpJaqzC+eQevAYE4sjqnt62HhJ1HPcFhfMTO3fjHyySyuwCL
ftJXXSkW9dqW0gh/hfKA6sOmg93bLh8vgy/StU+r7NAbuKW9WghmPN7hOKsVdzDN
VIEyESSKwMavSxFqr2Lv6bWF/9QrkPFkajRxlHS/L+p1TgOZmaqIJBgLVqO4IrnD
r6zjPF9GPQHZ+qkylHyQ5EWjoIF41PCsMI4HdSQhnlD6Ph3Yd+1VKIHDpJwIvYir
pdLzwMaBZRK6aVBZ/1xBX41VfRBD/PVfl7ki/xEAwzI3NqoqYjGxGAOkE6lqn+gz
zp+2npAdugn5q9tOYKaX0yoL4MHtNTeB/3K0t+Fgm3HHG3fYT4PDfpDnLc8KPwPW
0SiKQm4+5qG1oZlPc9Kxp7xkd/OFM9RlT1U8AU01XoTD1PMurDXaY/QDhj9sI6MT
a16rOrrgFbhm4c8kc39ItWHw3JWDbKRaa/XIdg5GCtZkhlRrAT9qPV1Zt8m3o31p
xrUrtHoPCrC0TlDzKCsYc328HG4dreu/2BHbuWp19p3r5275zTU3pV/aYjqOMsGS
Cr24mJb2ehcRCewmSdNnkU8OKBad7QZZWQ3P/dSF6dMdqY7Ts1VKOYeBIFvzd5Ef
cWHZ479Cc2Ytko9hr4LZXAM5vnoYYdpGgFzxXhQZ5z3OeK2vD2ndncqYlzNEWjOt
N8ePM6SERe1y+dEriSbAXKIvZTEttRAtLFIJ5m0KuTvQzRYLEKMBrchW43DToyVT
h5FOOK4bzsaD0mZdGFhza5DBaBJkIblH9XAjO/pXP3robio9QivV72P5fmICd6Q3
epiIFWT4ERB+0BaIdS+vXh53+h3/WsTSHH+qqJw0cppKsdJxBZRjonRNMaWko+VT
GN2z+Fncgkb912U+dfddC3RrkaeHqXTy4OHhXkzQxlQ7JKRWRyLuT5A3Z2LO4VKz
LFfVLD7crsojtTGw1rZloM6wfFvJtiCMNSghWIPKvqKjljCv7CuxQ8uuDFzSlncK
Jq+hBJtf3faP+fXDMM/JtBufP2Di8ZULoHcImgIgK7RLvrfgpJxMas4bHtKdBbl8
0Tu2TzcDexhAoiHzWrN/UB4Id34VBom18KBz6ngGlpW+LFsbqyZoN0HkhJ3unA7F
OxY7PrOJCidJdW0jOQviT473HkTA1a2eyKigIufGFhlYBlaSejY9QjmigBqpcEuj
13OTUrT6ZWvGpRaRrK9s7/3PlBhUOK8VZAyPaAMiCnJwGt0mf/hGZtLbgD1YKHjN
XUL5nsh0J0orOgn8VZiZrHlxbxUgR/62GXert2VxsI3rYvuJ/XrhUfjiVhrcqBJd
G17HQLq0ysZB2TICboXMsHXBGqARV7ahvqpb1VgNGhtXS2Ebc9nDAa0vg8MM+AGz
o7/7dFiuo0JaWX7Ahuw8wB1krWhag2emu7lxsll16upX8xdBKv/qGd04Oy+9l1U5
h+6mKcPVJmHx7GGJPHMBgr0c6J2s29Fj3HSadj3RjOIBglJ1aRDAvB9eLqRI14cs
s8sxzHqHStCKhafz71eXS5LdMfkLA2SmvHI3V2r9ce/eU/wBAsw/MhesQSlFmoJ1
cgnTcf3XLnMvPYRkAlusFQpqPsL+3Wi5v5zZa0NBqnRTkcQAMLk1H0NAVY2vO0gI
iDIneEQ7VdmK9lCMqgP2zaMez0gX/otcnafOluNaLaLWzb6Fp0ziNVSGY48BGbe6
JUtrBYILBdjtGV3VBT2QCKGwM68+RhkGz9rbDZSbfOjK45GVutS3R3CbqMTnQ0JB
a2LHUb7KolNzYuFUNDUFc5qBhgB3pG8e2/IB04I8/kWj2TBhEM6sNUqoKlxD3cdx
GrqA8vtArG3ZjjORJ3F0dntgDOlEID7IfBZSBqA9LYzsnXV2/wzO5EWTMYvmg59T
jQsy5WYhJzgWrbTS2GIJojEBu3iHTx26bFXBi+3dnOZAiZWsGqcHC9oyKeTx3CkT
Ue7Iin3J3Efo8jbviREhsiHvKOXlZZmvU8sVlGcG8d/lROMqSaa/lYIoFs39Me6X
ej2gdIZTTUYzUY2TJT1oY/kYvY8WLhcEfdKTKM97/wnbLGwTqHRZ47gX1m5LjRaY
/4f1k7z76IZsNRF/XJy8HSbrQEgFJnUSpmVnbcZjs6FBszc8uugyXEyK3UoeqpS5
3aoKMhKh+WK1+2BqW0Y9mt1r8Y1CFwQfqp+9Vyo4AMHbnum+E1LidiWFpDbrpETt
Wo864q51vj9w/2xbjpq2USMbHqBPRCY77cSpcH0DSF1G/6hg/UkhsL5O6ad8ZWid
AEYDECbL8dekVby5BjuNXjDevDz/Fw42NEtuleByBYLoKA2LHf9ndfpNsrbCebce
Gu8CqqN2AZQ9lDGT0qjxv3mkWhrRpt2ttXrj8cvZVKH2yS38Ggr2SuUZfNPLeki+
bjoOCzUs7A/8af4UWx5jy2cTLQjxUd+Z2GLl4FxDYOLFgYJQ0KHJiRTRhNBNSCFc
NfSZ8tWljNfaBaplng7XMHtnF3tadmaU9Vz+ZUlHq9gB2TcFsVy36CGjG/n2gxe/
H+C8+NhRwm1psdHtKV0690CwvSoL5D2VaKqGivKCchS0EdwX3BAnsvZe3r2f4iVN
14SjyZ9kgDrTqQoyK1jleL50q5KiqkY5+Ta4ghj+xgXYgQLCy7BK7mm8mJ3ZN9re
t5iJxsWNq4l+87LQA3/dWXrOqQw3F7p/ck/BbEO/0DNRT5YLfdrv1vicRjNqtjub
upssqPBxsxVIoUY5Kz837PsxceiwMKuSgLH6n0PG5lPd+yhWnS2F10OCR/oAoVDN
kmPzSOAnZ59wPdCCwKLa0yumvFsCwWD5BLs3y4eFE2yDYs/nVbTOYczjuL9pjPz+
TJjWuZZacveN8J8J8Mmiy13M6G105oi2BNwXkedNCqkxWz4yrX6kB4kDvuQX5mR3
X+ooCYpNlgGcZJ+8Jlt0mm7VlcR6CkH2klLlpfurxnOEsHZioaEcWrsWcuB3kEaH
HHIsIqomHAHUNA1ytK95MrDHW3HPCEUBaDndEbnKU6yAzryK48uKBPxI01v2kmJo
W85nPyzH1vFX+BBlAt1jniLJVwCbgLsA3wp8Z8G4dgots2bjVhj3VEAkUNByNDk4
1XV2rnwiZtorqdJyLrgTVBuqWaVCkiXNjZeG1cScycPBoUYS2htbxI4QN1zUpo63
Ff85OjUVMoBDVbYIbebdHbhdXQ85yVixq2f4LVCuq3RsaC9QAWHtX6bQzOquAn3e
famg/UGhkPTQr9nB410/O6WB1m4nCs0LFEST2bdSPBaOCxPUrQP0XHCZlxNKYw1+
Emj9S9XwE2OJCLFHF4K3iR4DKtmTDYlzNwD6Ht3rYqdkMZvtQBCUiKYnMLTf5t0B
PV/T3sfq3hovCYw8nq521AyrcwXmxQaGKC2AKPFJfooG99ZQd4/TSqd+xN5mbCwq
Xx0FVzD2pku73Oth3QFmUFH6jAZjZEEVn1b2wzcA2OXTC5ic1R6mzVX7WDvY02EH
+XYIUnF47CjQh9Q7yloH/hHrD4VeA0Gk8Im1xXiUkuyflKgt9y4uJAiwaZEl0eOo
mxcrgfINuPoyERDyMkqGCuEG2EZMXYAfonx2olxWsv9j+1TIV7/gCp5Lm/cK2fcx
DpxkWKgLSNrn58e1xH2iF7qXYm/UT1eY576keIIpqVYa/dkFwAIdj3U/T38mQzok
KX7hlmt7lceU27NnALwtPDjuaGbD3TiLFJWOaQdKB2O+qkrzBeCmzgXYkrKFSuVp
XL3j5RK31bb3zKj0kLXqJAWBRjhEfUv+8etVYZOt35b10ENFnFxRXb7UKr3uiPEq
1YTb/JnCkWEfjNBH7mj638ZshSvdeQyod0UvZX5pA6XMpo4OobhUKRyRLeCKvEGl
xOaKXy935BZ7BevEpmKt3lUslOzVCn+a6dc2eRMYsSuKRou3QJCU0QCCIWOWizWY
HqbLMgkd8nhXxjLCC9or6C+bsCfQmHhDInhmvCYwXkB5ESAt8JkxT9JxodthVSNs
2+jOyNNZqxD/OQFjr14LRsp40y+f5UuytZqnc4Ghf+FxI6P9uSM5mvq+OAjl6gtK
1EwcSeHJBGPcjyT2qT40F1GzCvYlEeV4KEDkQzXnHSHpspRb2MCN533cahLkkr6+
CR1XtyCcZUp89CIIZ9H3dqMHf60TnW7yqid2Isd7N8iTWCE/CSA6iEEIJzUK0onI
ezZVfk1spPS0TmIPw0ZHFIGFhq8OK3JpTiHABOTfTMHz1iHDJ++ZxtsEkshmx0dL
meQWFpNlSAh2HKLKtECy3gs+nK5sDNSo18yExsQeuWQ1Yv0H9m3/2gc2IhRA5K1Q
z5HzGr5NJL+AHCL8esFHY/k8IIbWjrMpKL+aROGd9Qkw/gy2OevZ9yWTo4R0gZ+D
TpvXKvRr5E9VkAggXoYZdm+caTSLlzsfpeW8q4XufiQNI13KtzQKLeTH/EMhqesB
mO0Ob0J9Lp50bm6J5UjMkeEKgZwrVmvj3SVPrbA3tuwfRLLydEOrjfKHdToB7jW4
5cg1mc6aEDwIryuma5LEFX+8N6iej/eSe8mv9zdd3I/LA56ByQJDtE5kOUL5kEo7
MpuaMRZpxnMAdTwn4vwGSwkDi3r/E4Sp6OnmIPZVI1N2a4l0cFHERT6Fn+0Vh8Pb
CJ7xxc0n4x7CSWnjtAC/392g7N0bwD1DKuMPGLimejNqR+mTl+HO4cnE0M9N/oVt
udM2hQcS4K2vg9CinBzndhPp9ZXrCtNGNOIBkNoZFL9tj/2cE1wXwsT5gV8iv6FG
iJNoBFZt8AaT5B0jRzN1h4/ldLVpVlih3mvFBFAgrz32jo2AJXZquD871HRxGPgR
Sno30czgzpdu/4aLEGukvQsoXwCDF6G2EuhpbyLOz4NwkZE4A8+XaRQyO82qN9bP
7qrsvlahvZjyNPxo2V06OjAyOI/ESjMRlsJkuhSCkJzDS8o4FAIQGnspmBqpcAXz
Iqfed+pt0udbasnWKe13+O7Wbd16sp79iz5rhokhyBHvYF9fOQZTnHaBRWK8hXpc
T339JeutV5kb9RovAHd0eLwaBQn2iS09Hn1S6tUYO++jzuK+GwO7igzVQJ8bYcCV
PwBAGm0GVWPtVNGIlKVY/tCLyFPxlOwPsJTt8w4GzqOc6PP+FCsbA/aJuldHpwA8
0CkJrGNI0iqEq7PhEBvxtWsXKBcJ73ExPDGD8NFVckjMIq9GC7s+Q67Gnmfj3uiX
PNtuChqU53AD+Hm5HVDx9QW2J7QNXKT8dEizv0GD2HYnqaFQYrIlpV9u/yS3v/iZ
t4wXh/VcQv3+ZsMczTm2GgFlds8yflxPICPJ9IJTKnpttBfBWrHoHVLJQSBokwK1
jxRwn4PhBjzqqer9TU6IISYt5QsH3FPBYFDneRM3HdU0ILl2EjDOZH79Tt48Irga
7VmU2rxVyhKBPOq2WAfKQ6TvbFaidPQBv/0CKrc8l2hW+QRMUzYxPhmW8abcWnnG
xFpSdvMJ0fPUqlLUlVcaBulQh+4/cEQs0wkQqHRd2fnv2RiIYNWQloAb7BIkRL/B
AgU1bvon4fbT1AP5KDpvFOt+1z+WE3u6+DgyHBXFif+OsevhkaXaIP13z56io3um
xVrOKBzKc1EQuw1xikWsOnrhKrAZJ0V6Hp+ckCt86RT3BDk/V9fZdigjlXyfVZg2
a2Hr1w98B0d1AHZ5UPW4ZPed+ThoM/roqHpZPjyJaYPlUqZ2NQLm79nifGFOTqaU
rdnuVef5dqxRstHnVId81K2awGhP+e0onYR11rPYBU2eetZF1W6az/gD7RmxYAUE
2Znm2+xgwRL7XE3aCE3yBnWYnY7n9qE52Vk+OHp/4XTsY7Tcxflxh7YpysUYynBr
sMRdeobStzF5SNK4pQbscAsdymo9y+Rt4zj/22jwSasUXA/aoHntwOlfXNFbuSZU
74h2priaPNUPmENkECGYwpQrBsxPIE2thUPQ7bTKdj/o0fmIo5XUC/c3Qbgf/WFu
89f7Uyz81reCdMbrO8tzfN/F0+MczRYJUdm+4RMQR5MpYx3h6KohjowIT07wM+PQ
Ide5capGB49Qa3bcbzx0/L6OamC/2JI+uMR9rXZt8ShgIHjy39IFW3BYVLTh7bMX
n68HSImEUF9vdEF9VM5W0Jv3/dIwuaVg52PjTDRoHO4o0+eHVMekg6J5gEBerPF5
RJCjCva4kChruin7M3B5YBQ0sNcustm5SgbLRRrEO9xo0WPkNrRf4nhuUAxBRCUE
y4FYO1kmANVvJ+y/xxva366Dv99+V1w/uO6MMRJjY9XuLQeZZJMCCToqOqU+Mwck
CD+l8qzmzZ9zjJRUxr8propiw7C3Vj3fy1MwIpeEzEDKN9LcK3YuFT8cHy35sU6R
3l0UWdWB71bhjqyPWZNylcAE79JMKWdhb5voYIiiBuX7uFNCWa28hpn7nG6qEFZX
qFyLvqAVJGZALrFN1Mz05I884yhKMHyGhabXm2rHcZsrdQclPhH2HNZVOsYTNQhL
tHMljrxPT4XNsLfPJP6f7K/2e6M2TnyA1lizCuD98lEUWxfu66bR/jYabe1/0DH1
eWLIyfni1QG+l5RePot46tVFhZzKd4rP7zJOBnVKJ94PlffCDIzbk8gHgHWs5RMT
2qMthDDfV1hMdQ10Ye/fKwQ3ZvBeNzq10mAce4nyc+2ijoXqJ51o2WSgaDHus+Ul
GaSD7gLzFjRo8jGP3jc/GQGaxQpEfcBXW5SqxgLLeHv37+EGlnHCP2ZjQiIJGDQI
GjgPytgdiXE/NPPoKKajq/G4TnaJ3QgsqTYUh2KqaN3HQdz3dV+6PvPcG+ZyT33g
raT3/ORX1enOblHavNKwQ+iJ3Ftdnkad0SX4OP4b1NlC+sCfwG/UrL8sMl6pgGQ4
4j9TAaJPhrpXRDenh4braEtBcwgD9azMNbqzizn3OeaFGp3DnZV565KrE84JSL+x
DNwudLq/3eRVTgUffvQQwiRbyZKjw6H6vPznPyxPVMaLyZP/nhrxzrrjMfVTXNI1
aUnsF6NUnyEezgZ7JSqmsBYYFG+8isftV+V6Qcb059DQXEa1CO4+Px9ofOffNqr1
IqOk2MiNy582i26Wt5VjkV+FQtoQUtMurr8NTTH4v5Kes8sPPuNxMsM1UKHqeMgB
oHFjzCizXxvWaZNpa9dNZICwZuAcNcA/fczgkFOSCZjjIo97c9oi/MPIdHNplSjO
pxWBG8DBiEapPv60dgSdK1+UCc5HvKrHobRrNWSycYwBvvqPp6C1+2Mo2vLk5Smc
D3GrJwYDh6pmT3WaFaZJrs7kpDEeapAbJ/j2zrD+0NT/SWxgHjqbVsF4V0fEb4ru
ma1StjCYsT7CO4Hq//J8Zxl8R/3DiOufY9hYa91tI7BmW7Ljoxd+FD6A7V3ykWz7
wZBmqFYjztOdwR1b7Dfiz4RcMcPqgR0xRmJq6A1Iv4/am95WpV3aQuQ+kVk41iG7
PKHUb8nKReMoDHy+N9FjoAv3gG/KVHSIRvGMIMZNdqAUf/FgQ41/7JPtE7P2FMR6
nVB2QRpjy57pRAFjt6MTtagTc//iatFar8hIAcA86kw7I+i8bUrdeCzxKaHpIr79
4EzsVZsQVtVqtaSML3pmvPwsllFqZ4AjrsP0oOhf1PfiaxqmQ38lSlxtNJzVXYdW
Ner2OiKq2pqxy7qGpQrxTLubId+d5e/cjc6bDDxaG7JiJqQc+llKMYx69w+ZvUR2
YNOkRNRnlfhR5pSFw66HAGREgr4mTcYupu+2uUFi4zhe1lDtmTDiAP/A5+a1o9gN
zGpUvYrE1s9FwzoBmQoZexOufSn2hmve33Po6cJKYYgB/ffADH+vazqqkz1TijvC
4dhxl70Y99bxmHNviZG4OqWRcK15m4KmkJA1PKHbBfaLn7YeiVS2d2aORuWVJYTj
brRh0zkngA0NUOGSUYjlWoJ+Xph801w0r+pYLKZ/a2+xTGp3HWSr1pDyyCr9a5Pa
R3wGN2bWfpcLHirvunC0SrjtNYiApfBFngHO5z210RwshVoIoVGH61Of/RlsTUKV
7nFFKaEuMQZGntOFt1OAGdtg8jUcvyJb+3pkxbex2wndcJiTewHV3dw/yiYGWkCO
bIiE6cU0jJc4M1Y2nj6EgPItZon83trl01aF87TQDAomb1Xt/OahUrsH3GkTVPKI
6jCeNqfz4HJQfmErquKd7KFn5vIK3U+Ayi1aBOt92MS47kK1hyhHPp0AM3wHEsAy
TfsS6mzRQSGXvz41KZtxLZC/rHoNfwqJEGq8n2AcvZPtINrvGZ169gTbz18BBWeX
ilPKxbsHzSDwS5USzW/H+V3bFJRwRNfTcqN82kR2bt3tIObP10d1Tc4hbvY+NCQh
hxLsarhMMMkFfqCl7X9t9V4e2C+FdKiCHdqZnbqnOucauOKUlm5fv4DA7F0jVWS4
U+N7FUCJPKvJpyIccJocVcLEYxHuCyxkDozY5CTSaAQHFMGQAfvzuBEnrgTOr5/m
2AQ7prw8Wgc8F4zBqDCPJNfKEyD4stn5P2eZbfA1zsq+u+7XzkPvLowgDF6vfKyv
Wth/y4MXg4hVNVIT5DJstEqxS20dt/Nh9GiW+AgCY7tZbEIU76w95JKi2XLanQq0
9BLpOTPmsN+el8xPlNRANWWD6b/3LoK8B4UcVhwp4yHEbkIjIyKR+hsyJX52JGoW
a4HhgaajhvkJgtqMNh3ciSqbOQdz3w4P6a+dQ9NcYolg9mWdVzLwxJaIyDXEfkyo
7NAq1nYshzwuOI3H3dALhXNAIi5XkKg5X515G/iqH2dZgc53k9LHgVLhcWbClhHX
PrEU/DwWjyqeH8X7u6TMn3ojwMSD80ej853v42EDa8cxCPx6AGuWSkApI8r1bPRU
9+WjTdZcwNVv7YzJUeCFaYTcMLa3hDMeQAygRApgjVehW/Uf9aNVpkTzzMMbxEnG
G5XNosJJf3cME8yF0D5Dp+465a1qmapaQOYIyKsA+Y3RzQlbVlirl56Ayrrcl3QH
4QFrOh3UaRy2XoQVUPPHICTWb27I3+QEmre+JTU77EM+LiEzoXDIUXKvfMJn4O7+
ML0nsqHSh5mAMlpg2nQlIvHgT0t1QRqI1QUhTVsvTyDSbNoC5mTxJLwLoQ3265ZZ
KwFE1rlTYgJz7Iq5sBh1nhcHLBBCVH8uKniPQajGnvoOTy3dSZZrkWIqRrKCpUma
P+asTnx0qm/LlaPt9Q9soNJEBduNBiTzWBUX1Z7HCIaQb6ddnu4veUUIziv5vYh2
jDYZSYMn7+ha13FO8AIlZ5+jyqi6jYsC7h2kKQM7GiOqbtQKKsxHPRq52wEkNuFo
VDdy3Uhs2LxPMsfgIKRHp/hO36va0G4Lqt74CRFHq1fm64SxcCGTwmgOwDpTmlvU
bGD3lXuM0K2p0autfcq0abfaTuLDo1tt1ZKixCFZJJ4lGD3l0CJRIS+kc09cSrIm
6lxoGbaJkHESNqwsRApJSoQF2f+Z6KnSxN4avQLyyx5SHRFiQ1XxvhvhuziKI4S5
k+bDb3p/eHI//FeJ1Tz2nXV1LD0qy6SXKNB7b9E9RwL1JQ+h55MDuFMRV0E0Kgow
A1zuo36abWkOatz5ArSt9E5f06Ep8Z9x39gJGoW7/Zswx8UosiNoJapa7eOhl4L7
1A/u5Py61ZFBFpGDNyGvYBfnLWNT0ZeRQVelkaFCkcBQMYWcYJO0OdrQOJBtSZF8
LwZPSTl6V/pGNntyxHphXSA1aGqmvXdPRHKdBaARYyYHvpxZmKBF5rAAD7UJrQe3
jN3/U5Fe00rI7p0NnsNNslHmFB73XzxZ9z+SUuua1QBYxcyBzrcemBfrwtzxCYAI
Y3VTtqY/xIhnTsMfObzMlVO7iaPwrkzltDVuQyOPd5O99cM8GYdkPWnz9ErVg/Op
nogJ+ILMUZoxzrsJ6VNcNWV7e4FBztd4lO0AL0bc3wRg51I9jQbnqjLiTpsblFYi
Xi7orqPjHuN/8Z66lqdZa+yu8Ai6n+y6J3FjX2Ar+bTr+eRgxKPTdv20g3zJc8TM
HoBbjBscMWtvUThWySYW8D4y85kUzDKar2S3Iihfu9eELUrQfhBgj7mdmmE2zBsD
+dvRkSoSq0wtbjSoZOOXoaDrwQ3WohG96HXw5UxEKcK33Pb7+OX2QqYVPfS7lOhp
zoeVBvlNleEXTmRSAHNzOZtKjBpIbbpzBOBKUnS1mrLLoY5B/pGIXKc7i5XrSmeZ
FRKm1Y+hJCyAsXicj2iDmBSmknsPa6JjpQ7Z5K6AZaNeueGCpHhHSA+F9cNuDxq5
7wLN/p4VZ/4PXJgSAXZPEk2li4lbDUIru/YHD7jjfLK7mf+++L9TANG5LbrXp/SH
9qNSOAm9M/T/KrDFr5Rn0+PPkC0l9tcA6jrksgmstXT027bGl3f+olVtwyg6icOt
7XhyspiJemxPJIACdNFRH9MUunGQiweMrQ73Md3+743GviQjeRZxxnh5x3tMlBNY
JjE5FKSO4CeWntrysTeHnwq78h29KUL721LDAcbBci6rSj2UiLdIxL6zIzUCDkAI
RnnuJNauXsx3QzPY8Fv3Vw80FsTn3oMYzOI1xF4LmoMZ5T+M/lmdyMyjmxXiMxC4
pj1wKqc5kQYsHLbYWbIscOMC8Xcr03I1+PHh2kKN2w+CajaswPKwnt6ZNqvi9K6A
zVjWv5LQIpt4DfBh7/E3yIVIB/G6goZmfGeDmrVjiGXyHrGhWNVgNEfmXV6PlAhO
3rzHabfLZ1fmHCbyjOzdn2Faih+EqL9duk1SFtTXgUEM/OH0kmuQ6lxGBRxKYPrT
PKdIATExfoXAJkFazQwDPJTiPcxtIQZtYKWKSzPQF88EtBgENZxLocN1riZtiC2C
FUby8CJ2Jw3C/2sP3pOlYBE3mQ8FouLP9DGr9nFD+MVWRML9cD+OBsSPysMj/dtW
thLfuZLxh5w+ufvoMhnZx9Ar65qatrY/yFRJ+7eK2ygdCXiHXaPFg3d6r/grHwGe
J9IzQY7qhkiZh2mi8wg22jSq2MUIlBI691A5O/CTwjLPUvaV34X0OFSueBBigwzc
y3BwmpsAJZC0SKq7d8AZ4E1ITy6pbYvb9aOq9m68RXYM64arcPuLIJBzqK/Lv9ra
XflHc35BFCH0ns5m+nllRYaeLTnvkxG7Y3VMKKIRNS27n5JTZAd5lbe0jii3TqhF
FS78eVj+CH9LUDRWrPuivUOjJ/iqN0L31W9mlee4VgT8+IbPhzllJ8fjKj/wG7z6
h06egG6wSkB9d8YWak3sbXHKxYXRMg3rK8e7/7OQdmuhIGfxg+rzWM19WJ9pBI0n
zrT3nfSrnlrnX+yQPh9HCXGtNRdVU4x8Sk6DNXIgVIXTpuSRqkoYKBJEpXAIKIWT
0JeaoUurN6aEqNqsrrdMd+c1z4DF5ts5xiBC/b3qBGRzrrs5wSaU1flA68O82haN
jmpe1Wj8dEY/Mj6PzZ/r6gvf0Ri5bWh2Z5kv54PLQWXrmwb8narUo4sDgCQAjoO3
sBmLPMkYPsAAHHEnqnDjJF+gNRDta2DE9aC3XN8lE1B4r6S+Bhj5H4eGrpAc5wF0
lyDQCkLfeVr5lUH24CTI5rlI64Bho1tu3gZGvvWG/gLk7UBLHMp7AQCEgkeqv/Lb
AWAwZ6cWtQYxGBwJej2KV7whyLh2b6xlNXDKYSlDOAGDGXWqw6AmNAdelwPm4rGX
MfF4DKw05iwWe/pqPDPk9JT+EyPjU6MQ/rkRhI/BGGiaLml0WwaljHg8+izfiuhf
/7Tv3QuLRYwKOrTizBV2RP6CYHx10jxPMqSrDaAUF5DeTmOtK5M/De4qxDJVqFkO
FgIdfJmJVfMvwFAzgVEFF+6BeiN2MVfbMcTlmLyCLeHvWiHgUg/B2ylA8rMplW4P
7ATXwUljRmqbTP0hdwuVX1LVBg6cTAfD5H7t3ZyOdJappKbAyBxX+iRZT9dT8y1Y
lBbWpxqZ3NIkqJLq49HDsa7mbwklW1aXyl1awklLagRLhB+GONvduQBhjUVmVpJf
k5H+ymJs+35HbMgI3ehx9uNcBNe+rQgU1puSgSY91CvIlVuEBeMNM+gSjJ3iM5Vg
PvzYlFalvZaeGI+WOVuerzBtEUYseIxqM+l84pQOZd3/Oub/FnKIow+jKbAXoPN8
xBKyCRcfNdfy9S9roIx0/awwhbyNTbAi5KscTXyIdREiYhGZnlGs4p+UoT8puJzR
wkhPKpj6/VF0bq5OeGlBr98DvGPUw7LWNJT8NpZgBDZMfcahEqHrewAcQsFUSmLs
U+39GsXt/hKUD3WuQ2i4dlyo4op3mUeYm6F95tD7OwHXZK5lI3wnaKCh4x9duW87
uCZtvLUA8W842YJovXib8SVoKFHy52yR0zqp4hpgWu5xie/J+2LTMPEUNGF3Lf31
T9EM0k+7DpusVLMC2tH1phU6IHj9emFrBnykTh2fjBl5bhyh+6+qd6OIxtzRqEFj
VdyAdNy65GAu0x1eHO9xduh/PRGAdBxlN+NEoFc15xGea8Kw4yfM4FPq/oMYDaw2
XoQEegQs/BVPsLayb/saBwxaFnHubFOqiLen+x3wI+qeJ4PyPtm3rBg6/8QsQaMG
csBpH11KGFZrbvnY5aWca/SVsR2OWkYJrW/kOtWCjeSz8STVXrQxPV1NY+8AXbcj
/NxAXTeBmYdIiar+AKkOwZuRqtrz3r8xtr9VycxNwO0+jh4ET2Q/DUfHyIQE/uhr
ouasorVFSnel9UcdB2F+vqt45ENAT5uNyKoQPVXgy2Z5xpwiVxZs4cS2efEzFFYM
Dr4m5RVQKY8y5QJDtvz0+qIAa0Um698DS6Kr0uLt7Mr0ZjP/mb6ZWJdL6/yyIm17
uAmE0sxpU2yjDQRQ4zREuHiseYgkiavh15uaPYYJWhRhE83sxh+mo2LLcIoBzeFH
9C7rLEdV/NSySkFlSMazy+avmX8wsI8Vhi3z4fPD/FoR1znp36oSSKspJ6ba3BPJ
9NMWgmieZAx4bFOmjPEnZw2s9EJ2h0HQ0Tn3OsUTok8O+U04D3FTmDB+scDUYynM
LMhb6WyNpkphNqx1J+3nnItpnnwxgrGL1ndDZFKQUHQyDJ7IJ365eiE9hLAYXe/G
D/EN0OZbVNXAV0e8C1bBdDw7mzkCrO//vW4NzUp5NSjBsyM4KMWXWS6VNKE2fBID
aDKYE1s+TgTwwYG9q4NCJckLQVCl7mGL+KffAsoKe8MuDHOp2O3Eh72imP5+Z7Mq
7F+OhNRGF6N/9gmP0uCSwDzJCVdUsngoOmsbviCFcMZZSXgMDN624Lg5PeMtEHuf
882Mk29OMCMdpKUbvWLhoePPz7bG08UmYDtHJ40LX/5s6PkoGOxRJkAlEXnAsOyK
bC0/x5cWzQYFu1diYFNWyeLMbQ+8nK3b4LoIGdH4T5KebOAkJAHfxToH1W+Rd2jv
wg/A47hEsMl1UHDz11FandJCJCXKPqJZ7xS2UWX77XFGzNK5chyHDO2OEFwwDWi/
qkWLvphlQo6d3nNv6B07Dd8ecS0Bm57DCLMPAOmm4u8xI7gCPyf7fN2T/5jQ1ArC
i/RNZNHuqzFK8o+bJv+91HZzuCr85rWDRPWomlpBrTW2pxFdqYwL34gnTrcLZVo4
Dhhpe6vw8xqmKFE3PTYgsJo8+Fy72Blif/2bTsWD3WTUaRT/bB5NvdhFQIsgL5rT
xw3ef2nM398yrzscrGvXnom3MxZh49qb0VDs9scpIGGsRFpQlIGnMNwlJG7lT/Qr
JUW++rYhRWUTy5ofoBOf/FwY7yKtKatBkY3z5ybx6uxLy7S2boHmay9IFe7CNNvx
Aw23MNLhzQNeD8pzDeAxNEsNk4ctQ8J1t13DKCqcyWAIsq4dKlJ98eoXiX2HDr0T
zj+GYxu59BIdh1u5PrXkIvrfwjULAvt0yHB8ks5TeaFPy+boUk0xBVmgvEoNWcGO
1FOoVqhLKmGx350UGk6XYsGmv3IKSxeg0nkazXXAj3H6GxWtIujh0079m9iO9aZk
z/hEBf0Mp8UuZr3Me4M+p6XgvkBWVFZyC/P2WiB63AEBfK8rtqOePcj7FNAl/UjI
CagH0DN59y9H7pA0e01uQGHay7NM64JV+WEF29Ew0O0oAjjfclr4Rz1sUdKIYjGS
gb0WhPChjCJepmQSfeUFKyDlBGYmRoagXJWwvQVattDj8lpbMfEgot+KFHoTjxME
app4MR4KKb6wgmyHRLWKzTxcESyQZDMoV6/NaRtUsKeCbOj4kihHXtDZAb75OnS8
eaIEaKWL5DS+OR4bErJoRXXksNbmwRmIrVblr3WuBIIIwF1/FR/kaYakscG7r7G6
uSBEIdPPKQkmCvD8HKC80TD+g6PTnRTAFCXjZgoSKASrtAwK16mPCBepvlyHa9wQ
ui/wBhfUoPAJt8AdQSJzGLYVB/oavt40YKxhOCLMMBdW1RniH33lphzEEU82Besd
TIOAurymGZsVy7gA0+PYCOL6tvpYIl+wv7LWE7tQ8HJfd4cEWPNvafwuFASA1T+M
VJtaz62pyyM5Jd4ZZsFI7LbPQ8AyFKWDl4jjCu7PLBl7iUnO9zI98h20UM/fMsRG
3GZ7907cPWTNqC55snLLRydenIPGzekhGGjomBfOVp6yOBokQWRCcFGfaJ60aSIq
9LK+ZriuDqsp69oQzYNr37dicUYn8hXopHJ8u+mAOW6Ah8cw9nDy2V0kW7en2gmw
l+t71qkQ4aHbFWJ8GFNfINaej12cwJ6p5/WyD0XJQKZcAhDPMlMn2tcv43UAcRAl
OPXhPpLCw2WqlXhO1LY2eNuxnYOcrdVJ5zCE7Tf3pm0bLZ4/ib3J6PBFOepEdt4z
Ai1cJ3iilpynGjTYiO0IgKV+RT/Q+E69jM8eZek0U3YBV4mjYJzM9RPq02j+hMHX
uYvEX3bbZL3HU15w4TjKINR8Fs6u5ZO9H6l648HTfvsXUp1Fr3Jn0m9ESSexodaV
/WWdf26T5NU4+aIK00WvQejFIj41tFH537MombrL6BE08uw9qBIGP+7GKIWAQxZW
RYykZH/LubPJYtYMKYYTfKGNca5cCaXaBpeEtzGJlHpXQPWEuDshBSgpS1D/zRKV
h8wAB05JwQA/Ui9K4+dJjReHb4/XGJKFXS4CrPajGP0rvj+1KTzvf/6/8Dm4GA7l
1JgINOGXeTor0GQLIR5TPA2JVR9m6U6NOmURYmnAznkcUJd0IOSu8xMGBu5pwl3B
WgrO6HDPtGKcYf/7Hcg+de9DZply9G+UzJdJH5kymCWToV0/2fL8iYg4aPIz7MJB
8te6QfD87yLCNGFaKclnEENsQq0nwL5CylaSF2wVMhaois8rQMqIBCyF/JzZ5/Aa
VXWQaeEuiz4IhEddxXNVEKxDt1c2wDago7JvKB8bO/81EMBCdhEu439wDht3Itpg
Qd4jeHdTqCLj0TQ4Zl+JzbA62etvVZwkkGhMFSR3FuD3EnhTcKeXaaBEJk3AgpmB
cVXLDjgRLfiPjHrpDkPOhOYVvDOYC6+O1YUuX6b/06wcgrA2goRPXRP3MtyeXnST
xQvu6FFFWGqAmQIoPUijdiNOiCDMHBfIdZ7RBjnZbgdrBNfXNwh60rUFO9o4aSK+
tv9t6TfbbnqVg4R7zAZPH/rNG6nAYlhjO77KsDqLgVce2nNrpSrvNh/Z54vDwtYm
QE9YJ+nE7+0J6XDluKzlfPVs+C+7NG0xPbzJWS3qDEpPJxee76j0MXXJrhGhtAKg
iGo46IhfIKoAgEhPlNGfs+qcmPvJF24X3kkWSQ6n9oLzBuaaYmEuLPFZgwXyNwlz
pQujNVNd20s4e7qJ+qT68Q0PkmQxP8UZsC47zY0V27A6MvC0z8wUMsElTzDVL3BU
A0F2+GAlwgiC12tfDBE3kF/7oVCas4HUkeKrNi6frnmV9dnpUTwckTnsBJYdFlCi
E9a4HuCIe+HrpQmpebzujcmjR9S89Lc3z5Qe8j5cou8s6RctBogklhwn4b6lcUIV
rz9KZGIb4QVn1Mv3lXIJed9M5NBcmtjIB/DYYzhsbn8yNVZmt/EjvHk3plcQEFzM
vv1aQgUFhh3Pu3YaAKBMCep9KR7k4rTocIqQV9wC5Jys5jQ6+EEy1lcHPzOQgyMU
F+sMszFx4xg3a9489qxnfSSjzDZKXEXiLpaOV6Hh+MdPQtX2hzvt3nZ+AjIc5Ijl
Mphzq3b/otx1wRHiYihRd5g7y4L2h99hO4G7D58uwg9xcRTSUUZfGNiApY6XKfUz
uWyGpAYV+mB7YdFQoDHttHq1vH1lkiNzBN2JabFQ80JNu3GgFre9vQUgfpywMQR4
plTosKZLqvSf/UDd3RcCqKSEO2qF/sqJpVJUez0wp6Zp6Zm968MOaSqq99J04Wqf
AA9Ozk2ZC+Sry8lH0lVoN6Bck0gew+2g9YCl5U4heRjDtYvedh/s549hGFCBJYMW
KBHCXm5KdeYhg9pefMvnJmQMn6rxM1EzUWUAmGBPdFCdvpK3IxtUN2JSNGKPWjaU
/GVoRT40Y2LADjzbdlCVwqn+n+TmxDNb6I+Rsea0pcyvT3PZnoPfzU6w8TSYXWb4
J3TomWuMFrrerOVg8rGmaejTLlCXo7InAlAr7Z+Fd45C7L+8+ggQiwF2oebeElHD
Yq24rsV3vsvyI7jZlgWf355j6FMVjG2ZQ/S2iDg8P754m14mhs7NiHFu7AkMQQGG
lODDRMBlrx4KP7gSPdl5TObR8PPBfdmG97AIorSJcQ641ej8M8i6xIgyVPP6+soR
fDv4d8GwC+ts67uXBh1ZCrgv9DU2NkVY2qdknpV4NUhL0LI4LvJawpoD6k5yonF/
OklRaRzwilv/fvgTeK0V75CyNCOFpku35U2u8mww9WBtwtrmIucfByUumgNzqTa2
5U95BAHVyhJmleuZ/I7O0AKCrd5OFDYlOnKOmxh6/jK4GP/FUK3E+Bn2z7tdvVNF
a8vxzslmjk+3DFujE4YTH2YaX5oxkfkt3uLnQNb7RRTf327V451v35XFGV7RDIPO
zcayBMN6+qEzHSaehAhh0FWkGgVBu+daf/NaC977p7oN0ZiJVDakRaEz0oOaFvWH
/H2yQTYo4abMx9jxopAhf5Tj3ptG+QuceNLeUN5qQc6WGKMY+/huuOOh43Lnhgkw
OHBo6nS9hj1HFpuntbbHd4ZcwZuV2YRGEtaEsk670GcWn0VCHtlBY/9geUUmtrZw
nL9FKTq8PSkOEDIQvcX0lDdqhbOMaS8OX31HsZJLjn73IzFgrARQI44AFlTFtuhQ
AVid/QJLIZPs0z5hciq+M1NknCvChSsyH2Tdd/cTyJrV1GHOkpwudRcksyxNTJ2p
t2To+tQK0BI2C69mbYkSzWNAh8DBwptIvlIU0+UHlSBQsc/B6j5Nkm/pGn8Nwp/p
zwlcAyNuHvSCIH3HIgC03FsRxHoAGidhcwsOIeOYn5yrcZ/avsw2My4Ex/HHOnMU
3XdKh7iAL+b1NDIOmw4FWeAjuLoyvHQOfTH6gWFWeuAOWGKIu5p3p2SXU1xlaq98
GMjummJDoo95pOs+I+pEBPd4hhEmdChKvXZNFub0c+yeC/in6yULwzEhV72X+ff0
aSMWSZ/+9yzzLYLbvKHb0za7UpKzeHfSNjLSKpSZtLOy3EUip9jQ0EhskQyBW54Q
/A0BsxSnNn1serDsIuc/DskZ/McOQl3aUL+TCHUkaYBgnsGhZJvpWVLEjKZe0UQb
7o2ZVbqPO2urlLQ0TlRSvy9mwJ9dKyvWafOrj/D/s7J0bc3GdQ5ITgo0Icj2H2nI
vZjUMRy9NFMX+taA7Z7sHi3pQUrpfZZ+eK9gFZ6kPO9VJnKRGvGcw0ODc2NN5t9m
vegUStws1YFuwZ6MOzzvWiNMlzpXA74ZeKEdW6Z0rdPijPx6xTu/w85mSKIr+Rzk
bLxGALNX5p02FsTMvG7a3JkMplOSETUHMd8ltmx3U0kiC9tNjcRmKa5NZwHeaT62
D3EKKLZDuM+9vGaHzQIo9KGPXfJihPcIhTX4mbwOe9jxzV6ziqiIJZbtdVtODnap
jrsDCh88ecrWMVjSzwytWbsnIAw0cYfW8vr4WdvMVf0Iu3syGR6YSi57po9e2PVO
X9nPmiU/xCkt2qgTj7Eu3vTwFnPQp/TQcQRqS/R1NXhJqkdbTEd4JvnrFBwPH4oC
1S42UnNSPCf3wsgRERd6Kh5PaYfZUHI1A342QRP0nVmIHGMKbLFxDKC1qPNOmNqK
h2Viy61Fm+yctbd9u0pYMPJiigyvYb4DJMzElpzyMfMEyjCtQVgKrX2HMUgj9olO
iGakb1yyzZItC/dZbs4AWI/G5Iuv/a8lC7OpZMXY9uBwr7igpVguBJRcU+0gnuCv
4/VMsjs4ncBbnYOsHlWFEFoNIxdw2dde/JjsnWg6xcs3JZy4fk/CWEyXvy6wG+DP
czzI4mb4x+x7nq6/9UgHIzg5vDdIXiGnNhjlDHgXr7AH5Qyj4m62j5rYAMrW0oVw
M4nyZr4Awx/ati5ORZjbnx+5BAj+OCXDuesqECpaLyGNs9LNfOyCau/IFt/5Ruif
fsCn+QU1RFo3+uT9EfKFH1PCC25DU3uTBF2NrmJD9AddC3rSPvbVCamGeJatCwBK
mp5BhlJoC6QHAOlJM7ypTtSS2Z3cfBJpwmbZwohU2bxCK338G+NSvyDC2W5CpQaD
94YyxHXwhSSgO/l2HKpz/DHUqDO83c+XNUuDqC2OT3jWOVIYaGpqz9oIxSXximxP
yk1e33YGPyZ8bGo01aDhg0Mfp7VWDYmNjMUpE2j6W2FAWr4avKLq4KziSvRgQBxC
S8JCoJ14Tn9cqjU2kfWWNHv30Ctn6t5gkxxBUU8xWKGeg8Oc1qAe0gwOkVF3rwAk
wfeW6kzKHkZsoC6us+/fB7ZnKJ5MM50AxijjqxyvZfjppmE0MYzCCKhUqrj9rBMT
lG+WSP1U2hDmy87jd6ae9PFIkeQg+aEqySKwvIEDcPvS0VbGWPg1BEtu2F8mOgut
EvjA37II2nEeWaRY7XLiMw6M11fEId0ezkADfhRrr16lbQepw+puo3AChEBZ3mbP
mZDy+dG5T2LkHHbIrerd27LPrZOYCXbsyP9OwdXIdgFLXMSVa3zR7alL9qlOMVM+
eVuV0PgxK9tu0QHiOVjtRxcKIUMSi4RgID5u7SSrvj3JluSsMUOn1J1ED8kJzLlS
oTCcITJPDKXTKKD7o+oUEwnQp94gu+BOxQqc/656WXasbCs1ALpfmI1YSQyKjx6y
18+j9iNL0Y7MFQAF3iEwjiaK1T7jmWDfCmgpEt9+whURJ/qIIFzgMWg93NHLNxc9
CksXlNiWVi5gMh26kp/UFQMesPSTsodTfFtdhx2qzUBFCvZCJq5pO+0ite3kWZL3
umdwHozU53tQy/Hu5MW/gWAR9PkJMCddPBiuRyPWRk4x/uKb2x2af3czwqR+6FTL
i3LXTQw4i6ZtV0zev8+9LwjZXtUP/wHD4ynCoODJGS1QWWw16ialK24kmeCzWNj8
HeFgLcwy++6L7OtTWjlQrtMnRz1iNLJKRUv5PyJQzY/jhgDFSgO6ibNTjSNyHK2+
R16/odT7lAksd5iKHFJbMrxpZlhhMwSM9bMxoTP1MDnaFSW3MJXYSrCDgrvLbOzS
8VMuUnsQ98GbvTFZ+hZZ4BYNvBx0wXl4/kI2X3yOdY9aMndHp062gO9tPsCB2lk+
YjfdFXmSXjeiv5FhQDhGPYbZlcumXmBFdoFsClIBBR5RyVorvsNT9LWy36BKZ0rC
inx7mXPXrDU6kd1T4LrD44pEXocYGE33pH17vcTlUKOsVNnJq00sxVnbJlBgfNBc
jX3ZTx4vRN9yYLkpk/rl/85mnMkrmx679PrwA/x3GfCuTlmveLraFVJdZpF9vpST
i7dCWX2uvLHluCPRBcVjYZZ1ZTpl5NB+S8DSMzVVf+3SD40DorKIUTdisd7vTGiO
OXKoSI93WORea1q4pTAovDe5Aj0WCsSyba+b2RGTz7bro1VQ1jEljStne3T/M+5z
0Y3+w0ZL1Upu8s/xnPqfVVoMmgud1b0DWY4ZQffAJEoQeYyokE0+aDkmIHR2t8Zt
zXCCP5AgUFbj8Ia+17qtmBGnBQBdJR9uW/XOPpJfUk4gM/9KT9q6NVEBn616T/YW
p9PVt2gqHiFGPDYefEuOZIhjonv+dasFuUvwYMNTgmv8l75txDZKzQZJnrhTnNVO
c5Cr01J0LaXotY+w6cwUnO+YNU6jvU58a0F30Gmu4g+hhwBtIK+3z+hfTO7RUScK
tnuE2xbmcmQiI+NKMXJl8ek32V/+NBPTPqvGXCqOaLKSUp5evs7vZFHPlqWzdMeU
2UP+ad33TVDHNX9+qr3aPi5QV8ENVZYnnOmPXa2O81aoQqVyOwDCkRcr9QzC2tSy
+jANorFJvKwb2WKKrGJnVnxAPwugMhPMZ0H+nt0kFjR0VzdA6NJPUle/YsFFaSWv
JXwU+91jHL726hQ8OmR5ZmuAYmE5A6dThU7XSWtnp12eP3zNXWm3RJp/Hq3xr1wb
UUse7MnNVNqE6IhjVA6iqcnoumv6CUF6OqiCf3bzqTooxXSuMu0ZInRF9fQ6WwXG
3nXEAMQskJF/LhMh6DABM3D3tazNMR5HPkFLdX30q3puMZX/D2rcI6eB12Ez4zyZ
uKJGlpyjoQFMrYXy4ub3VF4f7C9jEbyh0d4uOpCgbcrbZuyMx2g2vZ/1c6wN0JXL
LQWeOAJrgYbZ7iW9D9awqCKFPqZ1rM9KJp3B3WUNLzfxYmC8YIZbTL2uAgODwrsG
sCOeMlbpQxOrYHI0QXAsv1VGaD2ET1+tFJS5hEiAn05UmPccGOXR42y5LjRjnS6v
fEYHfK8w52T8nHYGiQDXMm7Z7+FQuDrhfZFkVeDuRjsmev/Ws2xQu3FE5wer3sdh
YNcIR5AWaZi7Npmo30KAiXg2s0TaxIKCQgeqA/VkJsb+y2B1d692UenrxhfmLIkh
4cPPIisp8rWqKG22h1g4NNXRDE5Lg+/zEdBNYOXk/nyh0KYMhnqX3hqiCIHMIHWi
zJOflFD9g/kD50v4Cs/WY/Dy6ThYlE7xdJGy1W7gv9WII/PashPrn9mD00+QqEb4
z0ZC71+zHvBwzAyjQWavHbBHZOEzPRVkTjC496FKlcv1J0BkJW2ktQ7MolnkqlqS
tFF4rMpeJgSEaRqXdmhb1m8qYH5F3FhKiUI4d4T72K+GWPf8rL17qLNnfA1ZFQWa
tLW2ua5p/L/lsWo9BW2pl8Sa+ku9XhycZotcwrY9VfPEj4ZzfFdVhewrB9uf3wR8
cfTKnWeJvbBA0CoJxFAKQKWT9/XsDielCWVrueI7VqkPdpRUtTSwmRDTvlfheXP5
J/JgVSAA9jlNIzBD31tCivzqk97iE4Xofn3hl724CLjcYT4Azua3pV91wE2E/g9s
x5NdRVlpLBCuSLOft3KGFM3Pq/OfFDlxuKUzRsvkCvgYZ9C6z3fGG92Bg1EA9Ds9
lzxmCaqqDyiiSBx+EXN1diwCRL/kC3aOsafwB+IIaBR+BamlS/5bxiVnIyCeRDqC
7aDbG1fiR+nq8GKKewmXarK8x9KJzgCFFDI33WLBo7J9wU/5eXKJKgiSgddh05UJ
mEVW6mpXv3o2j3NU0vFqx3zyS0/UiE6rzZ+JaFpoBWPPyRpDxKuOfICVVoHv9uHx
dXIizdIq6P3Hlm1493vyNIlNZzh9w/ismfBCjb/4jDVTHIs7U3STo6EVry6szrUO
dwO06dywfrnpqHEsbGHB97II6zNLR63RMndVrENUYY+0C9udGrc+ADwVbqVsBzH7
M93/bs/g6GbUZ8LqOnKObquDhUgtJiRiUCDa67zRf+g7xocfCfxwGO/hZTouRAMG
SZ9ZjhA2Ae2tnOUQRpj8ZIBSeHXPAWVzf5o6wa+6AF3sJad6MG+MHSFVWd0QCYAm
Vpy4+NuuM7n2IwQwWSXeQbWitAbdUKJ+So7cj2XVWWnNLPNJ5Mloo/Y8Xayg/ioy
Yvr9zfSQGxS6+/SVcC2NxEH3z9lGSBBPZZHpeSP+bLpd6nWA+DWlJkp7v7DMyJvy
6iPlclQV5n7cxRN8Dd62LlIvxtD1gw5rQWLP2MgCfnnbIPZLil33yJ/g8uaOZDze
Ct6vBQnhWz8OxgXRiP4eMfc1vmbQCBJuynU0lwMzYR0sbQrXL9e6woxzvaN7mnVG
waIYKWEB28MPFcNBdmR7+SBlfofF7AzutGwSxCuQvQy3ST0FEoONUffO/I6EEqhF
oaS3t3VAluYeRXmyNIqzexM0nKr/bknSEn3DD29sKo++jO01CW4l9FjkwbQuiPs2
ZsL5lKxzEf7gWwqz0t/7KiFD19U0Pad5NDdcNE6786BZerE+mFKVLQ4CM2zC2J2p
UbeF06BrMmvdn3p0lFduZM1XvY1v/PXogQIV2y1/CF9gRO5laQF5q37DC35mn/XN
n/NYPKw5CHPWHA6NcyPdGdSG/s7qXVcn0pA8K/2Ke1gYZUqpF8iihXN3ooZrEl+w
kY8AJllgQh3MuZseZ79rl/2m6WZqoRpRq2zhrKmL4Zqk88yY909O/AEZEg49nr4V
DGhOxTG6QoOGEJcH0ZwanS5ELO7jtBXxkhHxeT9KBOUsAYF0oW6jOCzrnoyVDboT
ndzZ6LzW7V6eI2WJqP0IoJHaZgZ/Lem0BHAVJVFAQFYk6QnV6y8BgGX5+M2Tcy2x
AZB9+ISm3/OYV2Lx9Ut5e6dQrtn/O8mGszu+6VDJ6PaUzvADAzTFiPDGZ0QKdloZ
h3yLFoNcnJBImt1DTW+CTn4dWjeTu3UMB5G3TU8gjN9ZLW+4n85SihFu/rNIAxmp
S+qzzMDK4Eaxb+EbmaXjYKJjSzi5npXJ0CJH1bCeHZD7gaDuRoM2r3GDJNxKmAh8
pk9misvxgpbfeHibTyMh4jdiSF7QDmvVW1acfZnkUPLjlJVPrdBsEc3rs99aVS5U
68ivC39f1BkrKChQTnp6L0OGXZe75JwG+CX7xpjKeO4/XQHRoo57Vj8gECY0Xfy1
m0BJgD/725y/CalHn6e+mo/BM2AZIH7grbXdi4/4TIA6BKjkv2rXogZ/ggS2TmHR
`pragma protect end_protected
