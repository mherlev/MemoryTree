// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
`pragma protect begin_protected
`pragma protect author="Altera"
`pragma protect key_keyowner="VCS"
`pragma protect key_keyname="VCS001"
`pragma protect key_method="VCS003"
`pragma protect encoding=(enctype="uuencode",bytes=200         )
`pragma protect key_block
H+:"L;T];@KC\O]5555#L>)'3%!YQ><\C,?AM8YA\/,+:QPG3N_=%9@  
H,>7Q*=^M)'KVEI\K65[)G<SU;8/,7TU*0=570P@;S3(VC"&;Q&[)B   
H>I1CAR3._8H4:V-K_-V\3#CYT$+#.W.';N'!)96N@H6Q[\]74M$#Y0  
HO2^YP%0*:<>=4D'X6W?#*L= "O5]N-&%NKRU" "TQ2YD4ZTD>)5K#   
H)CTI>J[1Y-JAR<WH$A;K/BXF+=+C%?QRMN^0A3.I8P;B8Y<]BQJH+   
`pragma protect encoding=(enctype="uuencode",bytes=3712        )
`pragma protect data_method="aes128-cbc"
`pragma protect data_block
@RH?7,SYW,2I[!'-D"@WS#+.V?HM(3VS,I;D*5VF[054 
@A^K^68'3DW8F2X@:B+T1+W/I^WJ?P8<?#10Z 3@WH0\ 
@=R+:??WIK7(N#_B(5#^,$F^,.F/M7;<U#(^LO*<O6$8 
@XFJ(A)Q))]7Y#JYJ?'/5?$&PFG\G,8HFWN=#4YVHW)( 
@=-OLI\9RTZ:J9'4.7J3GX!XP#5'R](!Z2LY&;(#TYI  
@=L#4-V)C,-='R$7/9/,JG"Y[^O2OH\[AY9Q#YEY&<1< 
@_'KTU5/!P0C+J/,@,Z>RU"4;9XC=C\I)O9F'X]=7[N4 
@[=GVF\5YA^J05I7LW$Y*^;9(L*(W>5([/-7,ZEL'39H 
@PX4MG\C8RV\<4:K7IYM0-C5CY;;RYM9(\Z55<A"2HUD 
@3#3[DH2WG')3\E=LWQ!W^A.$&EGRO1_6.AX,BQP8-X$ 
@R"V\*]]31IV)[#N&=W/V>^!XTH/;O[^=!W5N2^5(V%< 
@/H5:R80L/$<I'$^DAO!"W;=/$(P=M@!M'?*9"\3XU<0 
@VY7_D_L?K8$?0_PJ?7 -COZ0G@V2&>I=<0K-<5094Y$ 
@%/(L&!\3 <"G\3-4THX]'G%=Z9Q3Q?3M!$\B NIX#TH 
@CU\JM>E'FYT:>,W2*HCJ%S>-P]19>(J=3)2Q*8<7L+( 
@@+_]GAW7C9AT?#_&KP&7XV/KSH;4(?3&P!B2.4_ 1?P 
@#1]7 6M;?3JZ:J^<&LD&>T?.(&DFX&!:BPN^]I4;I:, 
@%1D6/2+:1+.YP]WR,H+,>8Y(K01F=.:T:N#/9)P/1W8 
@\XKG07'*F9Q[6Q$KB':@0YN]I(R*O?O=;OO5K.2 \@8 
@;@8EW%T\O"2L((30FEB<Y&MUL6IX.)7FOQ*0W^ &3(( 
@E5Y27S[QE8&^NSE7DXW5("&@Z%)H%Q?4)IZ=IS"D3%$ 
@)\O-@<0HR6*6$W5N)BXZ)@'O35%:=U^V$K8#U%(<']P 
@[GQQY=94@,*C+VV#JD06@ADG>Q*7R;!0P3<R&W57JST 
@TEE5Y4L)"5?<\!:]</7^/)#X^T)M*"BXLRDBCLI,=YX 
@.3O=]\:X 6_D0GH *H6SF=N!F!LUA''?<,WL!(9L]9$ 
@%AI5YD\[A(H2,OSD&!I*ZZM"BJ&\V$$SXH:5$6X&7JD 
@!HF1]>MTE)D(Z3S*7*W5@ZS7]I*S.%JT*\%6YR1^[M< 
@\LK1U/3*J; DZZ0,N89*L.4V*QEWA5YTPQ8,/<D)*V$ 
@4ID[SLOW&\N8M79@O^W]3ZZGB8";!(/6[-N!P'-T8%L 
@&OI%?6$/4F=W@M$O>2@@0#T.?G_[)]^YM73M)3I+SO@ 
@2'24T)K@S%$UR\L<6(V1&M.)0?6M"K>!BMI%8)50H3( 
@682BZ,'BJF'P6(*F^U/A56**'M!)3_:Y7(.!=CYN@U4 
@1[[2!T4/Q"*>CQWYW^@HV*Z.S0V(.9<=[Y_^.?QC?$H 
@LX3N )R3#XC_@98Z9V_BP)H$5'\Z= .\3.O><A#N<-( 
@IJ6ZQSUQL5W9,I*07TZ*7'-%1C7F3@48U:XNJ14:ZTT 
@70QTF<%5X8C"$UV11X8Q_A;"A,S$N%@A >TVAM;*FLX 
@(K9H=M?1L]5O]%5,AUQ*3%Y&HA?%-K(C4$.#^6H]X3@ 
@SOS00 ]TJ/O.=F[L?K$^L.3P9T*LZ]%@E<7[K&?J=<0 
@IBHVN+R[&X@Y*HH5]*]K4W!$.\D;F;#5Q6O@[@_9ZB4 
@WLV518)D$=7**<_#<>B?]I FY)_#U##DH:4,9N0&5X@ 
@OLIAH.GPAQEAYC[-/@AFA8*W:9)PV7R7X"@_"MNSIR< 
@ZM> L* 48%6G)GR;3UD[7Q> UBKTVV\G1"1B&:&&>>P 
@'3$@'"3)[E*BX 6_[+6:FD0SR\?S)">>(9_1/X=CL(H 
@CNDP:KK\9I.K1QR[6H-$#4)O'*OMNR*?8 9TFV9$==D 
@Z2U2X%2PC*%W#-J#^6&F]IPI2SRQTQ/V*SLP$!2D?3  
@"NM7$!?:2;G=R!IGSB4_&*\F+/"C//*AU:T&UXM I6  
@JU#0C2X0/XKF9,R.DK8XU#2I"QTX75$R!]A@KG?=J_< 
@76R-CL[06_VJUT[&@8+T&^GVTA8<C&QL U/ (F-=\1D 
@FW_XG+Y=.&4,6EJNC2)/$9X3=FC? $(UH6:<)@U9VW4 
@+^28A@@,9YH;SVJ]R- IB)4<,N*4&']DR/>> F_Y"F< 
@7@0)72 Y'9W.T+U#6,''NR 0HJ8 F<QS$O.RTS')K.( 
@!>+G@:#27K1;8\<;%59\ASE\:_P5_<+*Q:ZX_)+3G"H 
@]9P_5'N>4^<#*43_$:6N,7? Q8P5G\D^=7:+*9)2BT( 
@CH(D?E$;;FWDQ:B?%?%_BC'7TIZL&\^.+,\;I;F W'L 
@9Z,/NBQ2^<&+[3=MH&N&CM,WPL(RNRC4(2V4_F4,?\X 
@,(V\>-@QF*-(L^Q"V%802<-5-UR57KIF(Q4>GNA@S 4 
@44!WM@%OSQX#C8M)F^R!(*!]ONQ_3SZ.,]"75[%+XM$ 
@?G\("P$M+KN:<:B\\WN'GJ?@G> G[<RP!,3NXF9MO7$ 
@EW&IBY4&JO)>UR1<&""2!X<)K;=.K920RF?KRGQAS2D 
@6V9>8_8F1:>[IL2"G6]=@+)J[I-]&MN%<5O!U6C/ N8 
@ 'MQ+"=K!QRI@S*385%L6D;/F,MV6!B]"$"^Y0D)T D 
@JWSSZ"K!KC5Y27^VRR,%1+_S4N@5]P[I:>DG<742E2, 
@:;A_23Z7E,PQ@\O%GY&M8422LJ\#>2_Z4DF#,CHNKAT 
@Z-GIP>8BVI&%Y350E%AX%UP#K+@8K25K8YIP*DS!PN  
@Z\1K\#,:2S"L8XG<84U.6G(CZ?*7Y]]9K1J(<X1I3H( 
@J/TFA>;B$>;:QS7'W%N#R><9C4XK80;Q[D%)ODEV4A, 
@@NR(&8,813 BFVNG]C3"(-)DP\L9^24C("[YC/++6VH 
@:QZ8#]PH@+@Z0F( ,83S!G^PYW'<B=T")I% #%*P2G8 
@IED]<S<@^PMJ"^<K\Z=*01XYEK>R/68%; Q$FT<1FE4 
@8.,.3Z&,Z,+[H"0/"D1_YHE*3:<)+O!FL]^R,1/7UH\ 
@Q?&EEG"ZXVT5L/[J([A;0;/HD(J!*JZ:199B N3)_.4 
@3LM@=/%QPN]"=3JQ*K/G[F)^9M\)\C(>9#3<+D%4(S< 
@KF"!T;FUW#'J3ZI7D0CRSQC2YTL]J&D2:KE?T#'N4MH 
@W[B7P9*%7I*101T'^@@-<#^M'&M4QA!<M"?A@;1QM-L 
@TI &)W"%^9,R\I[&@@N0H7RYKMLHX W,2O&*A.I615( 
@9?)]MD ZEDC]'A TRHA+I_]A#G%HOWU;/K.6J!3KV6$ 
@;K%"!DH$IB>8 3_)(1)-?&)O9[RG_9:TUU5V,];?W8L 
@J?2N#.1^_!^$OF]G^0/:5Q!GA#;2)IECUUT\OXB0<R4 
@VW>'.X4[+/NZ'U6JVS9"Q?(G9ZE:*8;T#?)HC'L1PX@ 
@,C-J#;9,'0S)(V.?S+/K0:ZYV-LZ>8WS+)EQ\J^A^1X 
@I1QM23VAH+^ XB :IOS1G]M1GZIQD1PZ1D3DI5XG?2@ 
@G#K1&F]G6C->'\5U%Q*(9ETGI%VB/6J4L._$_/P0K4H 
@>ZKT$,*KY(SO#UK!S:R#OX.Q0W'9[S?XR=!ALM'>U6< 
@G?RF=0DW=SQ"H 0:F](BN@_H^H#(EQIZK\XZ=*PL7B@ 
@Q:_3ZR*QVOWF"'I(N4N@.:"9&_H8^J_Z8E:OBOO<9X( 
@2743Q&)':1:IP'KW\3T&5I-MNC/R^YQMH6<E!X/VJK@ 
@B]Y:#]<4P'2J/I:E $"'ZCE_PL/SSZIX0<S7SFKCX$L 
@'GYJ2)-+;$0]J7M,3P3SD,7^NL5M7SWW#)CD$_>7**8 
@1^1?>.X<]199[5,2 &6JXY<#1#$_8G1(^/T)3D( G/0 
@J2N?Y.*KZ]7@9_8H/"]T8G5\KV 4VI/+TGX)FVYQ?4  
@@>Q_BN5TR$$0GVKP8+>=H:E0-^&S;RC6?_#VPL"789X 
@>Z 9#7P5I2*:[2BLGK4QDY+LG/=\X LQ@O'=W95=2)@ 
@9@?I$;X709EA,!+W/^B_>YFC5CS_3)O&BSHKZ%FQYS\ 
@<+*+R#/RX4HY,K*6LE8F,5W31F2Q_Z7\?>#/@DA[RMH 
@1B=G7!.M70MG-6I_D(8@QU@#2%Q)(]9\S7Q-RZH]68\ 
@LT[SHR-S:6SK\!<>XFRQ:P,>Q>'OX(?QC[17>CS[C_< 
@GB)&\(  KAF!?CPZM.U/:1W WU80B>R4>VX!*$+UX&H 
@I,YTTQ"KNQ>BA3JSDCVVN,*EG#]Q>0B9G+5.I4*A"0@ 
@>8]<&V6I^7GXH0ABE^YCO4$5G0-\"WZS6G?[FM('!X  
@#A'Q<F __"-3"[7.1ZIDJS;3%&(QIM/[>C:)Y:LRPJX 
@\+]0?@>OK_ <\'%E$RW.K>58X2ET"3.PE<'D&\:P-R@ 
@^)\G"!='$Q7:79BDMCD^G7.IFOA 8!@5\@2> 3=]XVH 
@P0\,# *3/1RSNK7E+4AT61H0T('4MUJ_.$*",-0<]!( 
@[X G?X,)/RB+B_;9A^QFAB]9MOIA'3U9)5-J"DL4D0\ 
@6#TX8");X!/S()+'"ZSKP$WBN%),:3VFUOVGQ*GAWYL 
@N#K*;AHMM@WCG1;!=5D,KICJ,4OE<&-,DIN7LG)! UP 
@[RCWHJ>$&_"3CD)27I)*^U)$B;C:+* @>@C80[[%P-$ 
@@F,OTA_NSY%%T90B_M8VU$T&6LX+!;5/RD\4T(*J<<X 
@=SP0U6*AX%J"L=U6795XV2[#)1I]PJP!Q(2TF/GU2O@ 
@9;'..D+^/0VDG4)FRZ'4R:=F21U<A0QS_GPECDZ+XG  
@9O>+WHXM[VE,*AIT$NCX("ET+%2N%NUL8"H9VB*)C>0 
@UQQY2!;AJ(2[V9W233VHX*/\V<=[";,D!Q[SV6!] "H 
@!70Z4;#L4</^%.4=MO:NBQAZ1$DNS8WCW26V"FT%J/8 
@C ,V<1_230PW  *VTIP/TT8>2WI^;DKBOLN<D8O.X4( 
@W6A6\K4$T7Q.2F64.V!.E/8C=G+([2!E.FV&U@3Z0(T 
0WT<A<8A*$NK 7-^3B?GQ70  
09.S3 KQ?;8-0,S!%S>?/%@  
`pragma protect end_protected
