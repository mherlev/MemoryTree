// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:47 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
f3D+GogmN5mgRhOKL3PQATvN3lNBBw0BYjEA+RCg14QiaG2doAFdortqliGiIBWG
EV4G+DAarY8o/04IPEIGcSW53iEzcCK3CkNsVbm3RF7l2CxGJp1etx6ZbEK6uWMP
eVk5YPRs8e9PESMfbHHuLCnqKCkSSXJiRO3AwwnXO1U=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13664)
MAT5OcEhj6Fv8PyFlzMy3cdJdhdtspH3jv9lreTF7V6GcFNUn4dCYHxDaRVlYuzs
SPPeh1tWCVzIokJ2D3qkXrZIJFTYBQuV2z9rty4jpVD7OOt9UuKSyoL12oTcJAfo
6vcMwsREB/TbRYDkzeeHz29n6lkzGzuwRQEEZswt4awkJ0+BSBxLhj/IpUUhU4eZ
hGOZr5QB5tXWMkr0K1mlXbWIzJCwAytadqNIVsm7s2R+PaBVSPSALe643adCvWL2
yNl8yCbmc3pOdXT8F/9c4MhO1HlECl0gS3cIjUTIh60pMSVtXQS7stnmcv5yto9q
JQmIneMliB6gq1gqmkFHqq3k7+PYMxzhtJIn2CHjMb3jQY8UaJZRlWdr/6wNluvm
EjnPfQDQ4aXOKTYBukMMpZbzUyY5+N+C2IejXtoyxEkcHAsjCubRthTd9g/r+6ba
E0kzNsU2lOGwYSpB5rZLiGRwb/S9TvK3dQhrNY1AjNg7o1k9vZ+zhGLU524reCSa
phsVApHVg2Axf/qOPHUPOHWo3X2Lr6a0ArssGLOI5j3bTrBAN+m0131tg1nKXp+k
XjwtSTYpE7n6r3BClM6Ht/SU59fABJR5zY5bUcvj7M5zhnWTPFhZPscX8Htox1qa
EgMCRtEmlCfHB5U4HyP2jOvxfmhm9HnFwKwpKIF7PHFdfg/6KQhIDaBcRGLnpEUO
/OGwezDy5KEBAl2cJK3o90nvkBXrQTCJ9n0rzlHI1/FRLQANkcBBfo/wwhdKSeX/
/9CHq//aHA5kPYsJlGAasdfUgA55Vuizwc9CsPCkT0ws/MH3iBUywhJEo88ln3LO
EqZvsMjfJLWvW5iDY7w0oop1oKuFE5zCQYfVyyt0uM6GTdOtnFhz2Wd+jaKQVUWS
CahszRkcx33tq4cILMH+BOlTpLPcjzB12GVyrGjm2V3FOQJAyd685eYOTgVBXo58
eRshSu7qJHhWVk0o95d9JCwAjPVbHM8s0lf25OpC3LJpjnYO0tXWGiZ6cVPsG5MS
InAn/V4QRGr2hMuw455XgqUey8skInP7pVLJ5ZS1P0tp3gAKy/w1kXoz2455fnqf
RRWWzI8+/TF8pFBWabrT8o//xMGFJ2KcRRONGPyEyIEiCyVLdajdCoAvhMKDu6rL
/USgciAkeGs/oEAVrZE5Hj2sBFaQv2ObFlKYozNj/dh1t2FhJVuIXf++oawOc4F5
9BpOMRySZc+HM9gb2u8D34xB+vXFCx7DYwzb+ms7w/LW/aa6jPM01hady6yHdtPD
lbJujcscnlRMCqdT/35arD0KDeq+lILcchnYdfw2R1bqSeFmPIsRKWLioi3BcfMB
/DLR9LZATY6zhL8GOqxvWqIUtzPRXbmiVXpeZ/2t1lPDCSqfTs5Tcrz3HRF4R6cr
r0gkVfaqlTd0DroXQET3MXwPLtJ1o2ObdnLRX88tZuxUIHl+gt7DGnGWvIklrR8f
VEzxmb4M60QqTxt2e2AOeS+Ty2WsgxXybIAD4j9jDLwfv7a3hqV2K7czscI84sBQ
UkRb6KKpqrlUu+trC05Kve/Dm/LP2BTZFmHhVo2KXtFNaEKDtW/9WGX/nHfpaGuI
opMjv1B0rCCizeoiu8PgedGAwWEVNlqRuJqA6ipYQBtwtufG6+H2ktmE+je5Fmjt
byzTSBNfEvcGdJDWPXibyzKTMs/32+Bmdr+cfLbC6YWZjcWiItVWj/86c9Y5jGsX
+mo/fii948A5UJA8bnOHj+7PWmYTM51vWBsr4Ut4n1AVbfoLOEV2Mt9Iz4LEGVnb
qZsskJ9lwNeeg1pHwK4hhSHZHWLUssZ7iLSUYvomApngZjYzA+UZGiAbjAyfA4BU
dyjH2M4w0QXap/3CVg8M0nd83YPh1WRsl4gqzFg1BBeH4IGwwJHFbzf8uUJwaBFp
TFZBOXsiJjk6nxNVBKBnNA8V9NkpTjPHQQ/J1CeeGqDEOKhhz02EloE7piKoch1e
Pj8ALiGnLgqtK2B8d1lFMbSPWRVPxbV5xwk2UIqe1PBRWDqxtGRfcnJNUxSi5lac
GY7z12g5xUN2KoaEBfOFIwgY0kThk2Xx3EDPGGFi9cfcs9pZmsEVpDYbugel5b2P
hVq0RMJEMuGxk62pMXBANBHnITpWSAqNpI2QUMezirooqTWyyI9oii7u2ep0Gmk8
kkdwixkqdF9OUTaklzF7UcrO4w8VFxaAxrggYdauGz7KB2jlaMqX9m74Re5Davh5
SSMzKJb71sVUVJzhER/tXKuCiv3SKLjb94VXJ8pS5LdXJL/GcXaFq2zRiB1krfOU
oK8WBrsT6bjYVCfB5YyHGs8Hd1l3mwRh6Jt/Apcm2TQHCafWPtHLBuIaXT3O6Lkz
wIn5FOo0AVRnAejGXxNXHNgEbkK1rGtmAv+P2jBYiUD8G9920US5m0RHJoWbbDYa
T7MiBqw2yusjJDvdHkbn6tX4Til68LPU+9xOPPqTl60virsrY2fcJgSA/RSl9Zit
BR+R6LakSXs8UnZiEnPbE7WN1TasvFrnmCmcb7aX4gkXHPridlrbnAX4hPQKfBZS
rJx3yN43jeMxk+a340z2YtHYJNcQCWFwdWMSfQmoG52p1QvLH9/WTw4mZ7wWHlcp
CXYjAx1QpNsDD39+BPNHBuNTkIfGjJv73BTE1dqai2BFrKO60rulzZ/gsf9OmWmF
G97SBzIaj4OCk8E/3bVGLIWSO+QZSUSZr0b1CRCve+iyqt33eMiXahcst/MfsB9a
yQeqLBwpBhm/BeI1QsBOjRhCUGB4YcSuJO7jbEWqnWzVxKU0DPNJYTDMwd48fOoO
2fQOlYBrTI7ZlsJhyl66pTtHWAjkGwJNzs7+Xcs1f/ajqgxXy27sfKROLteEuL/4
0d7QZeQMP6y2d3sMxa0hE1qjA90K3EQzLDxwHy6JEY/kMPcfnh0+ebVZZvtksdFY
kiAesNxqJpQrENNvbo8EMSBtDrrK28Arxi6gh2Za3CzTU5L48k/I0RSB8vUyC83W
8MZ7mG6IlkHrAr95pE87YH0IuisQFsGJomy8dX9gRV2tE2wKcXoEcTQuXDxJ5Nx0
NtrNWYuMPmIx2WHOAuOtcK3ZD2aF/dm5ZGEB5UAbwEU6rw8VBNb9vksuIrCDWtxz
j44+MQpP5D6QUi6cUZIlnqxWYm/E6n2S3mgBOBACo55e/5ka0UubVlf9Oh1Fi5ia
1B/GeQkt1hElG0c73NZxVg9W4tTCYkRT/EKOtxI1mtg2YV6XIehA6PokY4IjJH/o
kG0augGEepasB7UgHRAt/k8n/xeN7j7Z9QAD3wLAvr1v1zPna2PARDUlxYyDHyG5
KnmayVHv8vxQL9OX232dJ62CkbdJaYf28PE2YAaiWpIh42yRcCx0LLVG9h01VoPl
SR3aIwbNpBUQD39A2G6EA2kubgje5sj3p/GPc6pjb6bST2Fve47QGvwp2+RWoMM5
P3bES1eFjcsQmja7iX7pAvfhCbpZbykFj9nK+aSA61QfFUTJRaJm1EUBOQlYNPFI
qjXX4TcFagVgGAt5gkWCkvFosCSCFOpPilL88I7lKU0+YcH48UNk1+brPvVa82tF
UyWjUsobSL20gL1wLec1hj4e1vi8Za7X8CUfVeXPFPblU9yVitBWecTjQnuYMeE6
t1bm5VdijQYPcxCkwb3uUyB+o3HP/7OqW+XMIPJRq3O+yGfVW8tuAvLwRMuLpZXZ
8ypf/nbaLF0HY8BpXz+PVLF19tK1brvcFbuJUG7JgAUS7/+Lz6cCFDeBiCv5x7Pd
mp++oO/wA3Yiep+gxerkIIihXo5awOCUgL2ECpAwS4SLqI/i138uxN95Nc/JMycK
CM7bxs/2M+YyyWA0p4Qgdoc9zbOS9566fJAtRbE+OyffkqIfZL5yCFgthtuQMBo1
h7IPa5anD6paw8EyW5YYFaQ2Q63h0NQnsqHJooAs27cOR7LSRhaxeRHOg9yeGR8o
YI4ygfpIjrEEhOOIDbOvNo2uihl2/qNhFxGhK7IaNAspVatgN+Hmpcniplw1iffk
xfrQBnpD7AggC63SjbJRHE8Tlpto7NRhFBi1ZAi3Uq6OJ6AQIhKMvzh9UWYsFhHt
ThJtzFsszHfOrzW5SwN4kJSR9U2peDSMrLfW4KhXC8kP90iU3dxAIqt2BHRET53Y
R2YqRpVwheoHM7/Z5GZbVUFpTFBAcmTepkfIetiaJRPPfl0VCUmArOLeuZKuWziV
oCdc+DeQH2K+My1+x7IsY4LnRduqbDSDvbsGIhOZSvMU+t1Eilv4LoYH2Vmd8sMP
W3Orf53QsDqolW1YGyNlyBSEzvpJbpt+WxR+LMjUPikyijN6vZrQmFPcNOLYtyhi
zZGW2Ghkr45xowS1aZGNfgSpvC/uijNMEa7X+eBWp4SvJJgR6FO3qKbMMV9Li6M6
yBcFe/Kv9vkqrgkaSdfhDa5ttY8d3H6+F62hdUpPWCedw2qtbkQnnN3nGLdA7pEr
TgqTTnlxFdjeSoSwOpffR925SKxbsvT/4NrJX+VruLzBQJUfFZXcvDtNu9x7gaCE
QqpK64adHaOsoPUVRq2aVUNTCE3us2W99n+OVpVrCo5+fRuOsYrwpghayiZSnhue
/smlNjn/fV7Av/FpVnEHaB2g09ab+fGWduBYAYOmq665fbMHm7CdZDqRIJk9H9wn
PDjfC+N84M1SeVFcRGvyArLi5z43VnN80QO580bpTGAYheHYpYY1obCa6NDMo/8x
RxczqVk1E2Qscnm9sryLFc4gPuZWpuv9t3aoSI/63GpgkEwfdn9J+KhzLh+i/icI
ZuZibzNzk3DXRBVNauMFZ75ehqEoh5dTeRWOzN7cfmTCRKbVLdnBoxwUoypmbnHx
BaIQkGqi1OQulNpPizhVa23+Di4U+fGgBXnnirDcB4bq/uh1muV1BZ0wrPmi9wd0
IaBcgOYX8c2QdydD3GCJ3LP8/fa4I4EiYLWf06W219tb9yXbwQvfMCDGKE6eUIq1
NEJIx/jiB0tLW34s0Lw6elx+o63DMZefKWRMx2GOF42ohoxh8/aNYzk8ksGrNPR9
9ZurMg9Ff8HwZBnCGvVfpTmrvjtGvPdKr061aSh1vwrePaEiIgR3ekMHGdG8HKwe
x6IQkUsgpzsNEMDzAC2mPSFbA1K4dsglnmGhuNgfpkuZf4h8YsM+d2jdyRKlMIQ5
QLVeCkQIsPaOiK1+/MqOsKbui6G/86R2GhdtzVqNrSTOpIIQs3rl2AzQtG+GLsUa
rLSDUG6n+/Rmjvrd7bnipQ7twMo/y1GIOLGHiNRljkgzpWtL/CzBw1eMpHjicmea
5kPbfyICa0S27brvFHwJAOo4FhXunfqRKZg8/IjjCh8MbOHKJU5pjb2jR5XabkT/
4p63UOQLcdDcMG5r8p79b9CRpIAo71MW3SiPE/GaFlIZksmfCQU5aQkBmGa45B9S
TJU+do+QhCr+JvEH5AHUuWeL4irH1tGPlcKKJYAfTSxVT9tObhZJJabAs7fcwzlS
QMFzc7XBpH1Bp6cGA5GZCxMKiJy/wjSZVWHApuF4aFVZ826+unAcPUqFUKuAd5b5
LbySnovBK+KvRlOmOsufUoI+/ErRh7GEl0iKYnuoxR+O87mGgTvOU3HVBzhXf+mG
K16mxmEZU6mFUgHStIrt7nSNkMv+INLHMFLjkH+h0iPdFVyA6C2sE5Uv4TzGcvRR
wFv+M29bVq0fxXpumLBeBkm6MQURMQtkiJbjQ+uo8BtvcvnD7KXfcCyEYJhbcSRj
hm5C+/0wkFyM0yewoT+ph7/9XJsJ+CY+juHBN+5fWP7SPcrYFXb8KRbywFDhs5UV
/AGeTU44D2PbJrPlMYMaj6ozB20a5jwBc25mAtU5KwckbbtIOMp1ppEm91u2/xyB
i6iqVq63AfamLGPfUFWu8qeKcthV4ygAV0Dn3/GIK+PNYwTlpHJefZGOIel99BEm
puqeIGe63gLJwDici89uuCXMn3oVwA1VrkXD7FsKusBPOoo8jLiNFsEtIcD8dHRE
c3WbyRxF6G+W2kyEnFEb5RL3+kb6I/B6lLuNgEgQuHSR7pbIUZ/TLoPAvbDhMLBm
KHBOrnTJFkjxZlIKnZOS2PVofpfZyxbKZc2dfQVCksWP4eWB0eNq7/ayAxigHuRo
JskLN8zgnlqXt9PEXC9JSUZn8b6qGmLJB0Cp+AdBVidw2hYQPH26V2IyGzsKI1k8
ZJTGklliuq4HTy7xbcelj9pguI9/kGswXe2qTr1w/SSeEw7yFcIDvy4df/Rfr+b6
jDzsBqB9DNB1pCxLfa9cqjOA7YWhu0o+J//vE4oewL6elzdX9uq1DzAXYma6hRwr
xJljmgfCs5HQlytFWWeaQDu99jaRAYtJSX2yJ9p15TxXR/D2OFd6NZlaKk0R1DDe
Yq34MC6DF6EjDfxB5rtamRlEHhH0j58qOxOsEeYlTY6H6HlOBQnr+G9xT0ubeQL8
Qkl4dqbcx69Lj4TJBVDfvM26VLaFBVEMii19VZ2f2ZAJr7AUWXF54dhFbToI8eas
rxZjdPZocZx/lOdGI9lRFG0lpYmAjM7JDJDFpeJ/DfXY1v9M6fR5JZpZjUCLtC9S
+Xa2T4JcEKgMUjVTuaoOFO9PVM9xA53YG13ZSmjrb3YjqVEx7NOfMgLFG/1tlOwd
CYLIQ/dhSN4kNnIwp51SfzwPRIyfaLMTFLSB7Dfm81NNRQ1sbVRZD2KCrSHYBR+h
q4KAFXWyRwt+IVuN9ZgP+xt90VMRY3p0mItt+c5NIRsRsFS28hDU4rEZ3TTEf7YI
2HxjeZD2t8MtxDyjXXwRGQqQI15aCK9UZfRke8+IBKlY8CsTeSIMNckmfb1gVI7y
NNxoJO2hPtPgaqtIADknxXCbvJVsbFaBLR9qhkBqC/5Z2PDT2HG0lwDp+6lmS5ZN
s9CN1C8vdegtXV3G8+0B+zwRRO9eNMMSi0cdDigSaOctTDNXeKTByXCEmgouRIIi
/0Gz6ukJz+J0fxlskm6I5QyhoZRCWN/JIIwcIO1Owd5b03L6YVXLOhiqlhLSstXO
v9QKrceaYkiitfU3Y6jIe1KQJ9dJgJPsy8BBgYYdeZXH7wfhBzd8RBvWmF0Ug+Fs
gqZtlPRImNC+HIh6LjpWFIV1Oj8MGU9zof5rl/k3miL4lD5LIo8ipFLTp4DrLueh
uxBRUF8MWrYmQAVjL/s1XzKPk3H2Y34eYgUzCXuKdeBKLScHFhA+y0qZ2nxh5WSM
YKREbMuwIZO3O/lOfMepLd7eOquPKNBx2jpeEkk7wzpxekGboXczpIKTQbV7F5Z2
Dva0tQOrnxhN5m+gAdlD91hBAA1bBtR7vPm++RPtAbSvMW6siRM216q3V9ezisS+
G6XpcDv+FRcL6cJhM+OkVl3Ymliy6qmeengpJXLkY3Y67h5lLF0p2l5xv1LRvFCi
khFz3runy+bcC6V4OtICzlrLDhysWwgu7+NjtWEaTkIU0XO7WgtH0e6IUfjhmZo6
etjB7O59CseyF647phA98UEbSBPwWa/GFOIL0nRx78HXzuFezRbAMq3PLCmlKY9M
JsWzUvz11/3CG4uYgLDVF0IfQca4fNbWfT1KJvA2dux03zDS/NthNbx/F7XYuPQi
GxdCLK4QGERYAllSiovw75u0HvZyoDB62Ud36gELTCkTEo6VxtqozijamQOAAdea
dSD5OzFm6xEnqV26EIqCWHkQhF7eRedccssKw60j/NE8CjOLlVbo5RgMS1t5vUUr
06jQWsok54aghBKidA3FRL8A+fSAjQDbSBi9rduo1nAPI/yr8zMyX7oKVmQ3ZROA
8xHCHVYd8tJD2e2C9M3+B/SVvNhKrrXq0RcOAvlUdadLpLJlEGMbBuCduUXlRFDB
IlTyAPvjXHBeKxUhFUk02abhly6bld9M7P/0swexldEaW0wh+4jCA40nqbJwvYnB
KRH52g+jN6K20F3RdgN5oVYRoBkimZc1lbGMDJSjOsXSV0Ud9fzVmrfqsQmqke+y
yosT1osYH3HArvT35pMFMugV0z0LIJBoJprOQQIScTcQqmeeOFJP6HY8jXZ8b3kX
s9RirV6vur0J7YvjmkLKbfiotoAprP1sWeXf9hrMhwd6JxQhUi2Hiz/XuIwXz0Vn
nKLpw0HgNVB1T69FP67KC5dM3fvd4fLGXm14pwlktVWg6Z7TUnUpMqs2hx22SEFc
6EptM/Kz1xTqwAeV0VTh7XaHd06S2bOQ2eguPMgfBaGGl2g5pAjUNxm25m4Py9CZ
OFyzHJfphX8MoE7/2rW1qM406SrT6QLW1FZWt5V2RfX8QAmZHkbps1e/ZRfvdvwg
dJxPGpcBZ7FMvJD2LKD7UVXoOepDKkw69MQkxd8f2B3I3XvZylXxeQk55noEt2zO
4yEeu3wtKMR0bNOHFLRHmbglE9sy3PP2lWkJ7zrHt7xApURLWv7/ibe6D1anfCWW
VAVB9x2t76rrzb3MDPPyvlEfdKUhgKv3wvY0D5GO71QYI1QOxh+CoOaoiK8T5rKH
sjueJsT6R5x1Tefv5D4mbNqciBuaA+zmbx5ff4lioPcO73ckrRYcKUWkMcTVj/KK
yEYgecKXz0G76zG3Y+kVYF9wbr8j2uEnaOdxeiDDF4n5/df3+WSQMi99ptyk/Tg1
2vrLfA0abmeIovCBmnuGUqDhT6vYTnJ4JDjnlicLZboaO7mG/AKCjqf6B9jjiYR/
+6Tf6hBs8KqebKL/MNik63TMJM4x6XyRfgusKerunEM/R+TrKOndowP90kdL3NW5
y3rQXTKg4lsJhXLnQa5YGhoKA+LngVyHjByzhpd1vzLKP+W1/Q+uN5LkdIqA3Ws6
ZO8Mz83EMzgwpvgptQfqA5a4mxDPT4PfjZeNvZFNgyAX/BGq43TcSImOeRkBZn5Z
UDGjIdL3mRcfwTX8BRTeLTIMFL+SuvpdUTaPep+4ut6m87JtuvQ6ceaw8QtUZrpw
vPsI+DAekMERJntG+Fd35+e/OvGCNJTv5q5Ah7JPCI2OVEr+7IaFF0G2XOK7lhwg
z9OaDXiuLN6JtZ4t+JGdaRRswTAV8o0GFW2a8wBzGAjPCA+kIr4qx4oCHVQ8ZwDH
3wLbMTe5lBM0f5vKl8xIV26OVYmeRmLlW9QdUi6ArfIhlc/BX9D/ejUhqjAqaYRn
p5Y09cng14dQ81lqKK/zfIF8TdL3gCJmorjlM9wiT8IxeCsFlhYqPgLX+ZNeQX3j
IQsyFfYqFiyjHh1p8a6kVTOQEzN+hzoumz8iW53sROs6BoFBiaPuf1fTvHzbKVFQ
Aupb2VYBqqVsqUgFsbURzZVZQoT//9uzV/9/J2VioVocGYT7ZMTniL/8shluib37
yWx7bBgMfPNBYm33RIiy2PXkwozkAhw4zpYbsj9H9w7O8TpQN9ss0YUSrCf4x8+d
MluiAJh2b52keHEdcAcJISJx1CmUIh6KbZjPfO7QMP7kg9CErNNhQTpBhMPfQ9NW
EjYXwTQTIIpUmLEN9IpRECTpJMPIlllazadIgKuH0AssXNSr9EnE+qzNTP8/3lqI
NQMfgsr3s6VSPxU5Lbv5e4IS2byC1L9tOCfzqayH2mfDK6e0VT2gF8u/DoAC/6KD
vBXHNlpyG6mu6/jtRzQ/7YeS2Mmgg7nt2Ua4ySd4WHt1m/BfVF1B+0/BSzTFepEH
ZCwz3NIh9nbDV10TdxvSQcaghBdKyoDFyDhGlVtCN4YwFIV/KbDT9y+WeT/425o9
qIJgwuZvgQZSoctg2YasLcgwL5BTQrNuvb8MgBnnqjfBhj/abDiAzGbNx0ll6FvY
ZBPgyaSMWQghv8c4EGUU2slvoaLpCxXf1hdilCcisiTNoddjtRuNOd9HGgZ9oqel
Zxy7+RovYLmPkHwBnKuWWIoUvc2yqa6zAtXvfb4bprtk4OsBSLcwlIE+uIyyeqWD
XmFd7K/V6dZfnmB0iDiGTtM4Klyo/XmWoVe4DNqKrv1jwqYaTXJ9oG9o/LG5dh4H
t0NFvn1rboJS/6n9HJ3n44Y/mAe7FNY5byPrauJi+SdkE0y8kRaGW3IxnQ4tmpr6
pnfDm1FLqZRwebsZqLjIDt/oT09VseQtixML44FV8kPtcZk0WG8iEiI7TOR47YOL
rsLN+bl/4VQmooAmwY4giKhT5ASwn4hGrTw22XiAwytcfCDcyBNpplD3hoj2QPPA
iUX5kR2yUJFU0Aw5UJVwSrgVPUgN0IUJsA+fx9OOEpR/QViGdFtEwjyxzmosA2Gf
MMqBIn7YQCOFIqbO5SKQczwnD+267rbynUJpYkICpryGHYxg8V4BAJsN0MzRTDwB
mvc2iihkMNgHZ+DH504GAKP9k7d87F/gnQGsvdDGcmbUgwpw5LrkIiOCjhW4cSlL
cgokJqRlepiRCMgEv6kE6qr8UV0gZBhFCmQAwze1+5EHolFYFGEhz3xYBhOaPiSG
RKyqvNBQ3qoU94ZontDRI6KPE9TAhh0mSqi6uzUIlU8K9Wu4KskAzQkqVuW6ZM+u
aaXC8TGNiZ0KM2Gr5LLlac7A90SSjN+qiCbAGfIABN2h9f7U/lD2bhvWhTNvKIGP
4+6VX0pwRPcxxFiX9YkTIPS+XWfm/AZtvCxWpOVRzpPqdmH0b0E5yY04aFNejHJS
ydQZF8gHFh1zSk09P0fNa1HCkr3unWTCHXSovRgIGIrhkbSYbGziun62IgMRxKn2
bLQat5ZvZtu/jde9ndO4bp0YdgQLPZG2raiapQdN4C4m5/c6640uTj2RbyKj4e0W
Ycle6Mx0EWbnTroeguYDi1KjOZ3d2aoFW7zMoXBY0f25eNrlMDWnVe/iwMaEYtkR
bspu0O0Q3V6u/tKhB3TbJ969Xaxu2rggREIs0vIibWX2lr4ulDOW7kRuwm82PGdm
EIROZzoNwt3tp62bHB22PMzp6VeYFYFZh2vZykjQH1ghfOCAZy1joO/Og66tA1AF
Jjr3pmHIvl05/qmEYbpRTQQoFmxzXdvO7Z1DuT9iBelnahQ+vzeque4Yh6xuNCot
29wIIxFzuG0xAE7cCIuw+cAHvDTuJD5O2E2UjpZypANKoJ4Ex6mQAnBObX4w/ysu
JffVybPqrWvM39+GLx34QPCqPmMv3ydXf2N6H0OKDh+Rpf7CBr1U8eaFk0PdIJLG
nVOeZ7zGxm/m0q27BFLy3sCCVcCIquZskP+ipeNUPx0zAHVQm2YIsjxFE8o0Myrz
aXPTEKVu/jQquv7UokmbJ1RiS+LU2aTsh74I8P9DP6mmz1zUN/fquQqzY1cU/NvK
fyGD3g3t7lvtKxKqorWlOLxB+1y76BkL5jN/pC9tLeSuXZxacRhJ0+r0NPYGDTFe
f2cFpv6oVl1wUkjfWJzTh1s0zCW+e/jJNnuYYIoyvMOeNfLP+By7Dxn7jGKBIMEM
6sN5ms2MBxLQ83I+eNhzy7MGbzeysw28idadEvu8HFNzhK6KhjWKeG/zyvJgWWe0
ppAQSBbpCdRpr8/dAoCrmpJUu5uPrjj6IEFogTz6ryPD0jjfXkJIwdcf0I7FILvJ
cevVGlZ/02nYl13ZMpa+AkgeyElFGBwt4bxgdbXHjRlc6uZX+aIGd03Q1MkeP/LY
Kz1Mhyspj4P0a8q731DMjoHTAX06Q9sSuMkA78t1u1ov7qSdgt3WzrPmFm0rb7oP
glYWK3zjtN/1ryGcrnZ+/81szUy7NW3GmwoQY6EFXOaBu6QeshVy1G/MbYn2Y8YX
quXh1zZEOpvhmYKYMcDL9w4/gBFADRhVkxC6+K6XkWKAP18vWzjqK9UOwsyrn/Da
eZirSto1t6BP6sLt+RMhku03iSz/InxXNqsRnegunMtxDuXFGnecHOU+JAIAhtxZ
uxW2KQp+T6Y+ynEj0TCGPEeTUQK1/YiMNU5wKXgOKtj9I2UqrGfFFAI2eDsUQqyL
UFl8Roo/aClBG+rcJkNIoF06o4HAhfAZgQxkI/u3bFlvuK7Lv3abwnH6+XPqlJTr
dGEBxjr5PeslBbJlF5Zh1RGx3J3BKuUT4pwO4YQtoWZZBglk+XHAltXtzYBG9yGg
ojUSlcUeAuwjtsdlHZP1cRPTmw9VObXHhS7AQr3Z5eixqvhONUAaFDYRJljKtu1C
H2nn8UPPcnADhPtDmMlL1Kbp4JdNdBDmwoJqKWnIB3h8XnxEXOuLTM3zhwCcBgR3
78Gzg52SgHRC6GKt0WWzq8vfFI4cVwRyNXxdvZtLdQBXtWiSOQOjHbr17m8Hw6ZW
AZAhLFKAXDOyXvX9s6Cuv/dwlkIu35bkgYQmEQdvgi7fHfhE2iTvlL5cSlzIRASO
42zaXVj6AF3s7jhtEEuhiIiCWX0sHG13upOOKEwZFqPm93p378avbVPzFF9fGAVz
J5nnB8WbIECfe3/FyWHKwnkQUC7nuymlpslh3L7X7DDmk+XkqB8G7XlQdYRgC+1U
vj4aVjza6bftXJ+IBFm9e5ZLZVq6gjP+Td02aE5dDaCSXO5jUddfjdRxHxLaFaX8
Z9igFgGrbNbmCRq5xE+uwHRAGlnKFmBS4/1pv2tSxwDZxR9e0sP0aj40RuLoyLUI
FvY2s4LtzOwnA/69hu1mW4hk3AHKuXcQkfBl33zG/RCbLGwEbDc8py9dEzzq1Srn
SDZ/hesUx5BWiWk1zLOyDZD4JdtKJJLnoI4XQEI2lV/iw9l3kg/gwD4HgRiZxzA5
xeSSBwIAXVsypXnWNCYue6seoI279fn3U5xpPnlh9ropQkpf2zxfsrHgUPEq2kHj
9xSDQGZJ6RDogNuqrmQ3/sLYZ3oNZLwaXE9THW6nWXAAgEmq51/gOqqmT/r3Igw/
eg3c04YWpycYt1J75d+kvbe8X1hWlkuI6wBWXvY+e+ttDsViiyfPzRzb75kx95Dg
tBJXKxUldyACTb1rQFbsvxVPxZfDWOWB61MVRc2e+lNO12gx5LqPozYe0CNayaYA
tj5ubgtqij75uCQ+EGrhGy/yDS6+ECT/bz2kW7+2nUK7DrX0tclafQkN/HcOCJj5
zxsCMN/MI+FOD0b4KVxd/cAnd4tTDsQk/PcNmhOXHiG5B0rB6zDiuHCCZ01laZD5
0Xo8hBCz1WurxnJauuh56e2hITtEhofXlt3s51W6zUb4qT8QAho9IXhhzX1QJb7P
qqAscnjMYNXdiII2JCoiiH3Yy2dgZdhTTe/3MI2ZDIenHOdA9dg+QAuZLC9jlabz
1dh3UoCFaKNXFbsKixZHdOyNhgZq7JfCkwo9j2Z4Jpy6IfcbrT2sZ6iR6uwYVz/+
fHMjxpBDpMUAc68amIy/M5XVOmlwXVZ7/sjdvVHWarUDO53GRNM+SuEGUPkDJelR
F54BnZ7Vb5pyIAvU8gJg5xAvCFD6ssXYQMkTFrFd8hEXx653RX/qCCcfEDCUSCWS
YRBjDKtlaKCsP4pBEYGDnSfHoWWywxNBlQuARzybYoCRnyRWAFBgzhybOCr/T3PR
9bRPRhd29sJOlXPGS6aqPd7RchRmNBBkbYsB5peaHpqlgr3dPIBxsQDrmQYUKg6B
xrWWx8IPhutTspZv6ykZ3pLyG0zNNZbUJ5hIsvVZYPgbDrfojdnUZro6BuLjy1me
xxRauChtN4a4Fqrm1JPdFtTvP1TNYjXJHMeUOjehNTzLKUvu3tYjQAxKypB8xR7G
jMdRfrop6OZDwCf4Q7JRuHiQZvXsYeAkaDtjPAT5gUWGB6qgmYL0injeXFzQan1v
lRTIEhS34oMWQHsimogu7071tR4LLazz14QDclqpKuiNpVuy0JnGx7I6LzaqtFFJ
Xf629RAXeNor27MFS+nCFfWsD+c2ZItBjkYWnssXvbTcBR4XyZ8knDhCRu6+P08B
Fmva5d+m4WnsMeI54DUBwFwyzcq/6sU0G6KF7xSO9akkIVihPP/sv70vo6r0m/Ow
Ae0QnU+coOUXm9kTxx79T4nPqCoY81v/1sJVQyYdG3/ELFEgOxY3T8Gvq78+YiOK
ftizI14VN+lkRNGoI4NzA9cjbJ5IeO/g08lgEpkCaEHk4z6Idtf9mQSmOhcymCjd
tq1aj7u9jEq6J80cLlyboLA9mt4YTWcZEkAaZScfAcHW5IaDY0gCYTkIOlD+nJ+n
R+MtTPZUvuUcG54cJUAkmH/Qa0CZb6YXcI/OqEWL6lM2lzAPk0AES984CrMbB1Ld
y9O0NZhcP0daMOiNeLfbaRUvPpsUOdberY3jgR5EKducIjKXnvwH6qiwcSQ/vGb3
qyGi313yJF/x00/iZraFWRoyl8KNwmaAB8iM+G1RSM2SMh5F6P61w2BC/2KRA92w
x5QCZTze/YOWMhWRfbgG6AqfiKjHs7bHlt+sjwJXONqiEH/BURqgJtEzsODxMe9R
BRiekOXR8iGJg98JlA7Ffh8e6Ar+XhD5PT4LvniHSDrZPAC5hGu58wpkvsm/Z95q
1DyGp4rNBhwlawLlYQlQbQXuEJ1NhOZv6qLkb1NwxXIg2plOv7Thsr5laMjNfv6K
tv3C+LrRSFzeJE8Ps/UVtaDxCBESKuga2Hj3SBM68Diualgry3bPskB5RnNqNbKT
JYJ9L3wXny+o4HnJD8lbAAFjzh/lUwz2sZRzBFLAWWKUHH0zbzLDincaVR5WRnQH
HHPlZwZ1ogchR62ANG/yiDLVXt8bIN3aaui+nkgLuhIjH5YYg+q0ddhVQGA/ltum
Pu3Joa1pRC28VS1foZbba6zPlIsZDLLWGZiLjYavBXCZIrbndurjQihs8uDz2j79
7cxdRtcFbLMzfOA7TPz7JvE8jRrByiB7h34zKQFDnvblpq5IQqiGjywaYDzyb5nO
L5OLRif54w8Q5p45chSyMgERCfXRHlQdAuQUyjeHVpT3jyhNRqozVtIccjasBYKX
H+5rVvD9eUHzcZL8k88bJZLjcp1nGlICoRyyM3580zgJs4AzuXkcfcz8pSfZnXek
6H7AHRHbas4Ez9N3aWkb1U+8JeZ7KLC/AbzKqNMx66DKR2sqCH5yzIi5JPpesRss
kHbHu+Wc2xWgtyUKDkvNSusB739RJz2hucbvx/jrerwIcBrdWDAM1peXe3+PJ9Ni
njWe2rDnGcU0fgCzbg/dzpMJHBYMKj876WxNiH8SWiyrqHiF+wvEwNXFy28nzjpB
YZaeJwGAi2l5jc+tgLhAic/TgEQiRKDsVHQQiPjKIS7WRxzXNoWQM1mFfXAthyep
LRAjVR0Ftg6LrIatBKRY9FpTX5N+YoUV1xa7VuaZEfFX8PkyNxu+j+18gnA34iWZ
YguyDN2Ji5JzzdOYX4Bw/V/ctoOQV2grVFyBGeSXQELoPEoSGikBSl71UB6Mxdb2
h9ue3q7bnPq5Zv28qb/ltho+qn+8hPPcVuFL6QcQMgSqivjUwOzuUr3Gqo24OHwq
jmj3orTokiIhgDgae9KROcWUshtq0cu1bbnxrXrs1MxaFAR+43it58iqNPzpDqTj
DUCAIRG/BMuJwzbMF4i0cFb1nyHg3Gra1OlzSi9N5xh2NFwotB7eiAuzEtG3N0ag
j3kA6LO+P6LdykiJUusecskgoLNttCI0+Bj3JdC5cEx1r+ggLZDnQMFKVOVluNY6
LuniuunDeCuXUUtxGQQxRoGPPEFupfKWXo4QJs8jp89GxnsGY5Vp4Z9j7/hXyLgT
sDGZ7BANdYck+Ic6YYjvHkL4UKJ2Sym4Ag+LMy2uQeALZzc21hUQlT9TXKaYiEfR
QgWdbkhzj1Govmb8FHfys9ouLZWovzTCtq3ZDa2jogkfMZAIeuT9i/9o/lDXnRbc
IgEUxSj3wn7qi5t6+LFVm37Bpibulznh+MJDctvalUbdnaGFTehxjZpxsyVS+KG5
2QQ2NXmHRIUSpOH7+ErPQUn4Y3MMPHyR2gHKMlK2pR3ECGYbk3hhavSG9P/m8EYi
rANV4G+U1pp35K9llmojnAzACnTQvnBxEL4wmV2D4kexXoTaCAFNKlbRxgodKCb8
j6UMhZwyvBVO09dSa7Xeqx6tuiK3K6isM86TkIySAi+X5ylbRYLnatQI3OWMbSR3
mQwfKUxQzu0+SX5Kkq0/ptRYVlHqSaZeXj1zZdeRwJUwnv+wbib06RiJ+9BFtUwn
5ZgFvWZAHHQ+wQYzuIVCyMsmIY46DO/mYlz9uy93jIQhZ1qUdKyQLun1rexV6q4Q
qSYwSK8ALZ6YfTuy/zmBVFnIxAoK4hUUd9xSF0UUb0NT+lhMROGZDXbT4IZj+X/8
x6LLNxMHhYDif5PEIVfXaghYonKOOWqYyJudOC/SjjTTWesil7KTejNhIg0Zf0G6
QJ7qW+0CnojVSvMklYPIeCRGH1fz3PmnLHpwuEhEgO0YICQNI35l1xftPbNBW4C3
GcDM7z4YAPqZGavFNdiNLOVWLYEGjMgOC+OXJeQ6ealG6F+7s+FErlUhMB2uTRLs
t2cP5rpRYDhkolXrQdyJHZshNk2nlWaj6aGXVGLk353gFQonIMeRqy7zF8hFz2vV
vB+sI4/+Q7F6rJJ7lj+HKnPTm3iCDZluAUVsOhdEA90B4Q95RmSRkoDSxsd3nnjR
ThANmA0FNkZRL8HqLgubcKWu+9sq+tTwIF29JfNtFvKEsSfbyPFzKQAC3lTL5RIN
uWUl6QGP7KzgVCFdjJXGc69Xao2+89rZY8rsI7vlJDDQBBqIms9xK9CMyMxt4Dr8
+grw3lLhG7gVpokHkrffzqWLpw/0MN6pGkehhplo3ufL9qPtlyKcrHxvNKgam72D
LHRuzf+N1K5PdC7EjrAoAoakkBZjtrhw++8f8cxtqIaGW2TlIMMvWzbBVw5ZfT9e
GNy99kYMw7lzSKKWzC8P4YpHFG+x70GCTAuvx605UuUd92A+Czm9jjrf8Y8TwKlc
TU1dsjO27p+T6z3jasiNt2pAcl71r/l9/jrJd6ILpYgxKQhFzH22DKh9fsJDflJ5
csxJYCGCf17O5YdYkz5iN6tNk4Y+BHeMTGoRIMq7lV6Ye+0uS1gFoWM8+apos7gV
3H/qfpDVsDaJbYe7TX3x1REZUIlVdDlHN+hJFiWRRK76kpRsISF7sBFBct+UKtIY
5okHQ+jTh7tlTmKKh9Uby+qQ13XMGip5DPGn/LCkkJ3POqSqEZ9d3YoVMc9V/slT
gEzv95oWWRZ6rXAUxeakk/hGG7tC6Q75VtLR1QbCpkEnnRJf9T2MbvAn345qHSfS
jySu89GqrACIFVycolCqL3m5XDR9GwA4qHznqKq0uxU6KtT8Pab8Tc3ia+61k8sr
hcEwpodC/5Fr49RR/VzPCNP9DadJUC44QQ+u250F2tMITkAlqeq97fsZsY2SgkR3
4WdtewG+b0y1az8rpnIjwFI3cjbNVxH9bqYh0HL10fooEYf0gr1TeagvClfha1jg
MccxcM03cJDy8dFhR6r0l6lrz93C/XtkaszuE1D5LJWACaFW4LlJBSz9aQoeu+wd
ZaCoJqLPhQjXpy/+Fg9FkniHEcq+W0x9tSp7vQxfHVJm+IsAo6yfrvuApWwyHYT4
rw8jQv3ufzq8IVEINRJNntj40Uximmlp9HwpyR3w47crpDaJJ2ikzmQb5Se3ZcBm
GXImy1WqsU7fdckTw+pDNUUXeC7zxE1phSP6wtT9MQNp0GxkYTU9KSeAIfBss35z
tEEG2bGVzHbCe+QFeztcrUWJsveaAao/DMKEa7og4i5YpiwmrpVhLT4vfLQabx6h
lO92fa7okZgb+gUZa8B07lxX1MUJjZtBA8iIDq7UiX8h/T2OjFVhGC0LB0IiUqUi
nE532rXE59YfFzYP3coC/l6r4zjchVZTl0coM3IopX4QoAGOgOxF9x0Hbt5XCVmP
zRfyREngyHJ/U21kvkrnbMN9i33bqxzevbbYIhJuiQJYz+v0qTxZTfg5Wxdw9rww
ssB+tWu+OmD3A7Kd3iY6Q65yly3bc4zRszDjG0tOj8FmJFFKnUpf8UlJyWXa1KAH
32PfrWOYZ0ld4NnQzhjYl5ZGR5UymwGKJQRuFewCEBazGrgJ7gH3YXqYqUKQALzD
bIazcz9vDLXiyiLB8S5AMukF7FF8vS0OXX+zoLdb+YiVNGYedUr0mTy8GkGI/qvX
fdjusrfuxuoq+fNzXjc5oQbxJIIC24m2c8gYBzozTh1bf4L0BlGy8+bKa4menIUR
pwD6+YXppuQFN85fn5Uv0CFk13uWbjOAA0zLOjP4M6dihlaiclZfdFcgqXpEtUuc
aUnMYreoTQEtyote+gMW/S76dKUJkY16tkhxb3b5fxg=
`pragma protect end_protected
