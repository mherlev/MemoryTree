// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:54 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Ht1gKWJVFjvpUAlJo8dFhJ5Q7ql1hUgbrC1CeJIELE9QFj4ql5EZBbzXfm9uckXC
gXYmwr6RQOZg11rJgQwkA2SNjuwiZE2YilB1e09qvoWzA5AYdgU5Pfgg2RrUTEeY
XGsUuu16WTIoWoMZiF/VD3d689vcbq+kANrTyujAPas=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7424)
DDj3DOWGM9GVyIiW6muUJ8AD7Dh8YN1DlGXAKJ0+ZYcgXE7dHmOPztonux9rh5df
Z3kCDXxgMBhZHwA1YAfNGSC9MCcn5+WRWWCimdQ4NCDvs62XSWZI6x5tQES/uKu7
fF5tyS77QksS5FDdvxjw2qUuSaARfbuczH8vsmoGIucuzCjUTCtCMYSheq4sTPMq
rkUdeoKzZbKOe25XD8lKb4NNpIvyRGj20LcKwUdTaKJJLKNqXhRXupiL4Z1NDSEY
iMmpE2u4XbCGn0axFXmnt8z1XHH3U6Jp87amtbgJfvZSV989gIGxqpDlTmytxc/Y
TtyaMOx7qQAwgjVDuox6cePcVwXiQ2ZPeK/h7Pz3Eo4B04Pa9sNMCNuD92aLLjEa
gLcWvYmJgUUtWmkHo50VGNGmqMqIQUfbjXxKBFLNzBcfQbom6N6j34Ef4rvsQIua
7lN0cqzCQzuVhGPAn1Xs2w3EgMa2tZiq4pztx+3gv+WRCS5HTPMmg8VVSWaIK3qV
/ina0M+S9hGCzuQj/IV80PdAFEPZNeDt3bEOCSZ4i5R3F69Gz6DNOh9I4OwyAEnV
OnZiac7F8xCp7cT/dYgNYUxNmmzyOGGM9rIjwHDESSe45M8CPn1VXbDpKY/b20B8
DoW3sGALQR9N3ze7chBO8E/QClSfY9fzZ6CJzW/w8Nm0exQkitt+D+gvOO4YPeGU
NfEt1pc70fAkiEcDCwoAmsMODfmScNM2vhNASro47iQ81GFuzetApjairhab133j
x45NxcLXxhfcrg2jB+zBc02L+zcKtwcaGJnWnxkTOhALMJV0XNQTglC2boP1d7H9
L7vN86XNdO/WM8h7qiyqJwfB5zUDfUjKEIjALZGyfKIcpGFCzukH7j+TyQLEazjF
klDRCY7wUlz3rriTZ255ex9Sftus8ah4zGfK1nM/5k9BcccyglKhsN9efLmzl+2A
M8MwWB0rgxOpP7WP3tUNeSx05NjfEneiWDh0KuyAownIni3er2C2fLzWwMW9cqEF
03EpMcSStC0zOAEEx9Np/xMF1POYWGwYE9IkDdX58l+V3u2xO6ViRM/aGOHAzEt0
2hZdmgobsQOviHPHG4mzuyYhh3q5stYZ3Pglb8wkm7TUJvfvhxFfuPwd4apvwCWu
jqa51jWiZDo2NYeEjZcsnXjYHEsJya9Xk434Uq0cv49v7yBJgWXHgd2UHCsTYL1W
CnM/l6yz1nyY82VHkJr9w+E3LwIz0R+l5QfL9hugC8DQWflsohkylOfvfZ2J8f7L
hZXluJ/NND25cat/6a/m7Y59bLWk3DkEC/lP/pNmKuEnZqlk6cK/EuFSoNCM/cjf
HZwx5ztgT3U2UE7gngzRLGss9KYp/bDmBORXZIZV2VB0Nc2hIY/pV3YXTrroh7vM
23CiKwv2OWtdo3OGOq09D+KbDVXTikXlbEM6yx6E5De9XWmE10DFeOCmdIoNBB+Y
24tefkFYBdo/hXLBg60+TFRn41I/i3Us2WXYP05UjdhpeaE4nptkVj+8+8JTeLfp
NRO282faz6FEZsfxTgxkP+Koki1GFFpF2JovHKY23xyNMN9ZIJhnZXGthu0yYuVb
TLRko0PiqrqEZ0lR4/BBTuFymo7Ss6QZJTpwcOlOztLgafrYg4k90ZjYAxvPw729
RGxs4rdfuCj6rw4VUmgHHBZZc2uqEK4hvcm0n9gaFt5K39VnzZXDeCBFi+iwiHdr
T696kivg5w57QEylRad1dbFF+nxIC2CVF54IAUPSXfiUjLUflZVm8LkAkkCNkfSv
hDBgagPUieWuD93ZUiPRy0gzICVt01LXyQV/aOJ0Lxuc03ooUA642NYXkYWis48n
4zmxjqiYbuMmW6ZX8JaYA0li24J3pGYAQOU513VSAUTZjaY4+5S1FsZjtri+aJLm
BG5xLw/9b2Ma3jMWcTJfYrlkj8st+Eh2vdKtuFNTPu7I/cnXw5FpXqOMK9XGWjjT
/WO5gCUln2UQ9aOuW+pwdRPjyOrFwyhNa5PBnc//V7m9j6Mwz9BTfSig8EGxVUUf
arAHyf3kvZ/M73PbHFkIeFBcueNzZrn0mYuzh4QgOUjtOFKgbYj/78tgPjCceb6q
eA9j9JYREoH9cfN9CBPHdKDKaZfq1pYNks8FzhdZ1Rq8RvWYelIpGPAst9h+GOKA
aYtWcNCBW3Zncber3AZ6JxZ3TxOHK0xb6Stm8KQqyjAlPD5przWJmPeRRzdN7KWy
gWq04lbit16zmGt80rScTta8h5Soa0NZ88K0qZFM6SnLyWEyxJaYf1w2TLALIHUY
JQ79TCeR97jGj6LLw0K5Joih1Y+iQDL47jVK5DusBRnlMNyVAitNvYIlL/pgvlpx
t4WY71VXJP5MutINo5JpcOpj9c74CdHlyi53YhPsRBwKM8t+PT7vxa/jB/r6ZwKv
gU/+J5k2XpPme6JYDBa5UvCyWu+gsoPZIGkdrvyr41xtIScG7bAM11TnDwBLQXIk
b9iB3AUGTlV6lcxfahrusMm3S1SssMm0kg7sDcMrxZoYTThQii5cJEXcM1Y+GSYq
WZpJHRXgt+Ru5Um5+uODSSg/SYdLUYo8U84+mzyCVCbZ3rBFNPxyso16ntqvpBcJ
nhufrfkdHytY4A3ES9NKiyIckltH6nhYbobuL6La13C4NCcAPxbK+rEVps6nKKOY
Y1eD+CNH1a37aG4HiHlrelnWk6Ss3VeTO8bnFdg/QUr4EstRlrHIF7g/lp3up8hy
eI47KQmybyh0jhbSlDFE7AW5aAcpphorZGWYbNNOiH9/fRxEoTLkCKsPKoKAGllg
4mFs45bPrCui8kl/wSVKDj50/H9BBzXWO27VR9iEZCCZ9UOexNKVPCIR/ps2metE
HJvIGwrs0nvhxaNihgmJ8YnYNGqBtNrrEKyP+c0IXO1EVtcRQzAr1Og9Zpmr73/z
XHcAVBgOKb5anbT63OVnmXvtLlPiLtYpIYLQsoJIy3nqFE+jCvhPY/vfXbaz+B5N
151sjxQqxUtyvpyES/QP+D+aGDgDaFFUJwnvBaug9OpLwJWj5MRIKaTElInL7NFW
kdJ/7p02DwVeMEEQNz/eVl1rUyqvLa4r2lqnKXgDT9fpyYPCucpPBu/vAqNctOmo
od4mfdLHNCn3xiolCFmHJH6CQbNyJTOMwJsvB/DCe+cK+SbQipTpxFYcIsZuM+Ct
XzkzRXPigcyDSCkpzjIehSR9t04SF1FP+gmgnbNuySQjw9d5YT92k2yrjl0VL9Tu
nu2KPhb8naY2hwIuFAwHVNJudMuxKddSUx8lwSSj33zVkpwD4qEwIbLTTugA0iuu
R5sgvuL6SnXBdJS7I5zonyu+QWL/rB7ub8z9u/z9o9xwZYNJtR9Y3K66Ab+GfBv8
QLOFztZzbRfTDE4gw0/4jkEISUo1q20LRUuDqd++AGwYvs9n50pu/zOtSEFCVBfk
kOi0+K9BZOeBeX1lLjm4GTQ2b9SYIKiEy2IRTAxC8T+D5Cm5I2jwOJG+IeRnNZtf
2UcrNOq4pSJXEszAPj+9JADWmYGjjbTgyNJ2K1dJks5OIwTJstnGqWKoobgMGMZg
1xHnRHJq/qYRGFEq7xcfhftSrKxZE4UStp3FcOqrHJN2HAEkLkpoGy0Rho/wa1B2
qingIcLWN+W0yMbg/FY5GYmnEBsWAvhkKGJLFdDKeD9nQ1I9h9O4PzPUqmwAAKYT
Q+GikBCRHMosFOw/3uqSBH/LOVnLoywJqiRZBGtf+toqMgITy219fkjQ+dmX7H9j
0I2LOBIAx48DzdyKDkRipsBWEsUCeHLm+ukOGNfk71+8ADGUO9e/+rEcZmjVqggr
JfLDj9iqaY28lmgeiRycAx4FVbi/mP0qFm69MzB7OwRMg3dCk4agCGp42fGEcRF8
b+3fKC5b0mXYMzyHQC/qpT+/a3crU4OJe4LUgZs/onNo2BZTfc+mQT+w+Iaezji/
TcfRRXx4TNmUv0KRlFYg+G2Z58Y8k6M+cpBYYgIlvOcEAnY2yYdaKUesnOfxgFBJ
pJ5fpmyBPUJy6iNwSY2ibj33GDwWLMpNbK8vpMYBD9axUYh/cYiU7w1M/09AUGSP
FtPHIagME7iTJNCmHEfQ9zoOWewZbbWJp/3Ji9A89fibHEsrz4Sx2ijXm7Zt+sFn
CsNSMQgG+E+2hHJEP5aw5dlWkxo6w2Z1hWF3Ei3ep+oDMaEfG/McGqXLUkQAbc6e
KliHyG6+JV12EiDTUiFk2vTzhNrAlpQ7b628fCzwMZ/yrkoqUK93lyGlM10F3n/l
hez/s6uFhwjoV5zrwsLy105e8pq0ebPqwso+DUjv+A7nNWuvE5lBppuMSFPbOG7+
LD9USBW/jCmtw0VnsEPPSZDF30IELyKAuwC2780Vcoc+7OzVmwFxNoJsXAafszOI
mrFrdcduk3on3fPcBTSfBMjTr0DxBd4iB72amp+RaKK2Ei1axsS3kg15yTnJf63J
bfjkRnwkclHpvDsQp0Iwq5lQIttN2/AGsZdKafMre6n3Y67hTFnsq5UQv6RiBsM/
UOkeSYqMQKVQ5dWU+Bgt21oO0UFF8XkaeocsQSp+5Mo/PDro/g7UqzINUZ/nAQiC
5Z13jeQy1LT0o5sVFstTl0M03V39r78wrPW5Vu4FqczRCJVeM08tjiV2Fw5NyG3k
63z0rVVZuDpdlj/BTFqN4i7QqPXPw49pyIdJ/6+3pn5uKgGtKmBLkS931hhuvS5h
XBtnEXIheNvc2EN8BRzD7j9l6Co9jFlyqw+bpEp7RfOP9x7jUds5SfaS/Hcd0X71
d+ZnLwbBEEqQqAD8tAlAR13SV09uW4PwKcXAgiSdsM5pYZdsb4T2LhDzC2ea5cVK
w8jQE+99dbo4Xpi51Hv4tmC858/rokJ+Bpqo8BHiSa1isEgsnMkm8thlFe71DzKp
27VhCw8OQDamC0DLUTS8n4tSr5he9lMUu/sMm2584iVRD3H91ZbR+MMmgscEEosf
Bfq7Zt4zo/tM6PS1nLUb6wZK6igbM6MxLZ0HLAATK0rSUdhsDQfGMeyz/pfirRzB
rsQn0xudurUXDbIaFN3tC0YY5bYypBhIVFvh6M+3LDCMPi0wQ4EirzbpFP4FEoDg
mKt1UhM1YBH1JpAiIJfm+RsvS2AZbHpW9fq09nHrakTG4ToXpyjdAWmj0DWEIvC4
ptw598J4H0cNadn+mRcqYV4JfBB+Tgi+IB7BnKSOis6dt6pYd9mW7jjVWNvQXX/L
WNOnjP3Wr0m5U6qn02f4PoDO//nx93RYYFJTeKz+rskXcQ0rRoiYLG3BLk6Qtad5
ZqB1EISk4i5jCFG0zZ0DCGzeDBYIpA4WzKHns7fZi0wsp1+7UyOoceKa39MUZs/a
GUtyQFDzo03DPQIGQWnpFIqWBW0l4ioMwLsp96RLvq33hmkq3dvW6X/14bVfdFsk
yyrMSUlkwJibvArvvW1u1LnfaUOt5KO+6Qi7L6pNAiaPIVbycSDJZVV9Cjpd2p2i
wegdTD2WfIn1Reeww4ZZA/fXXyy84VXFEgoupklKdKJpyLlDDhRhSQw9lZAH4GQb
A/6WiRqVM+MQ7x7QZskj0UZHpF7klfbENYffq4YJJOwYKKux1L7O+7WtejZ0DrH7
jfIpolIk6qJDHUGezro/u1c9bBrkFPevhBgyo1pgBrwA0t+TcVUP4Yh/b/CbrDmR
aQcDdXF1HnfcmjdQgZMTr00AP1nkK+d5Tc8fJsWK3K81gfJsOQyiR5Mv9bOd24/1
1InZ7N8a1tbKglLXruf1aFvZ5GMhdZ1a7c4vG39zGZZMHJmFGzbFvAdj28usteXB
8t1l+dC1NNP+GW4XUTrJcv7XupfI+/N2Amqg11LF6rFHrKxfe6GlmkbpK4/46so8
gnhi8LFo4foS//UqnKnsp1mMw5nQ8Hs4z6i6SpKb+XDY0Kb2pUhVRLL9bKqB9alC
gE+Tf6OXg1rmM6WZBZBvgoB9tEIzb3EtgoWA0jjX9eqeJ0Pl7hOV7HgWzBiRLqzK
hok+1KkVc4f0bXezOIbGgDcfmi2HLdmhgGzYtEeEPhARwZB7Mn3bCmR5irmdRB6z
lH7sg9p9IMqQkNPgKti2yRnVaL64iWWSuLyLSkndWgqIM33stwILlP/oQQIypGK8
gu+kSZn/Ef9maMWqyxAphZCmujOSNEPXkt3wWIGNquod4ffiItNOu8lFaKOJOlpG
ewwMY/k3E/qVR/9oUKdkv7cJlwHY7hwiLyP/MV0gq0D1Z1WXV0PvI3OiZmbDCaTO
FLVb9Dq2Bs4YZQlXHZu/3Rnab65+SvHH9AlFoewVKnaNLVjEV5Qz/RfICeewJw0w
D0w5EIPMWKr0v56razUd9Svobl4m9g++8kCRcvuPu6zBI3tbaaBq0Up4cp4MVfDS
VQMulODJswORqvpbntka7bpuQ5VDuWE9bmKNV/IuQI4P7YRQUqUZGQwcC8orlfAg
qpUUCupiOX7llcxLb+VyyP4m/rUndoUSdX7quT6cudQVJ/GRu3DhYwAduuBkPVJF
qMlXGnDEO8TtwG2SrNHAYtJ3zQqO7oz3WJRZTYTK5G8FQzW3AnCHsIYWjq6Uuiwi
BqrZ9dV1bxR5Ajop+CbLbnsDuKtu0e61ddHlHd37iHteI/E+vfED3TUAa6Ld8pPP
X03h6cIT8WsMkVhly2aoBKkiUap3L4QYcU+D3oLT0Hpi0Y5i4cI0hA7I17F1MGKa
uWi4MG67hhlLj7dxMkiW/xOHaKilGDpbyI3VY0SQ9FpRlRLwfXcFO+smlrCpT29H
dZcFvSrtozsIZWKKxVyktuDYoS1rYqA5l81jQhf0gJDjX2ynolzShD0v5Q6uw7K4
K2pq3eDw6uY3CKRXVJz3TMb0cAQjgqwTOibSaWrz5yQ1AC7tnQ+t8xJiMK8uS2qv
UJ9V13ZX6Nh1prs02oSnMgFZAQu9m9oUmg/2wsPNMnLT0I/6cfbr6QYHmcVAihCs
rYNJ7grW3p7fR033j6jo2apwbu/iwAjAXGhNfIyM84eUJR5UY2I/VTdTmmasgbFY
WzhqzzFT5CMwkLkxe1ncel86UR8wo/U0ol+ijmxq8jSRepdA4NvTAbMWr9pcXSNP
IZTbyIS4orQotL03sjYAn0w0XadKlq1sObxyrLtK3/SL8hXyFewBkTEnkYcAlF+T
boMBrKHqZAJjwpXVazO4ivNa4D4tt07ACeEV2Xj2phbn1DBPPTgAuhp4BiFYkzur
EivH+iUqUOCH4PsfqIGiKyo1ULcNSsJ5YtKlaDZEfYSqEeH09wQCayFmpdoo2HBm
2ySK/OLMNAioIro0lkTmCUqs/Tw4L24rCE/aZtV3OgJejQN42UtYwqGhWqytskPh
N79Hgtkup2n0pmEwA0+XDLzRDCBbYmcbzlK6xi/FFY6ACvYX2IR+0YZuSJQ1U4mq
elIm9BDNzpe4Whph+dsE0MmMjPI3oycrq7Gd7K3v85ZrTQZuUgS0xNS/6ifWzFhP
66bWQunnN41ZRjZmIMoI3i16uXyX4u2d61Ciwi+S+gy0A1k9et4YwYs9bg5ccYwA
ZszaBcq0862kNucpOwU9LxAWGEKOqHbZ2NMSRf/cQEDlNTYFD/hOh2g6aX67vFNc
lF9b1Ekqj2NDYs7GoTAPZMexN7Ne4Q3Cbpi9JU38U2kHXhc+atxxSpwRFI8sjR8n
c0nPQLsDQZJM+3q4/px7wvgfM1p0o+VoZfd+dMSrKazUtF/E/IsQkR68LA55lc4L
zcaFH2aXrGG5UGBm9eFAKMmMdj1qMSEX5RkBz4D6JIUtzHxlvVGHLpkiS2yTmIh9
4m/kLoN5cfp9bUYQ75vwmPNAtMQWnIGrdSqF9kzHJea89KSNv61s5oi6a6cs11Vc
5X+tTFh1WiUvAWuSjGojocKpF5BNddm3itxr8K0kV0GgEZLISSm6Lh82glwo/SC+
w97EznEbsc3ABmmgGP0lnpj0ppgbqxdSZFOP28MVC7sKSnI0yLeLPH6RCbsuAWeA
bHhIxsC1QiGoS/PfB7zdrqeXlMxTuLDNHIfHSCqU3UGFNmPZMKDUgdh6CP56RzR3
PvbVvZRyFXCcWrMJXX559FjXkzBFRGszBuiAGkGfMYKbzDpUvuhWhrIcfZcjLbdF
ygoCwawBNNGL3Tbxp1KZbD9PeqcR1+tHbL3+nLItD1SEvRt89+/F2bktA/DqDPoX
+tBm9cD+F/eSUOuG4Qui8sWbyMbqZMADNFpD6rHp5cIB9Ev8Ods1fWRwyd3mB/uE
pQYnefDx1aMnR6IVjhFNtrwcSh/6NMdZxRd6w2thep/mfvJW0ZLLmFR12SWEHFXs
VYiQvJnSDeFCpZI7w9+QIHZZDqvl8285yXADSos5LGn6ivmDnOrPSpBfzrKB+aax
/oS4P0d+CFHbOykuCVOJZXQXvtF3id/Bhnuh0U9fk4+6QL1k2QsMJfPiMsqXbjPi
6+i0r0m2lke8TOwWlRW4JuS3cU4Y2rMU8gRizB57O0allLMiK8LxxSlO4hqsdNB0
JrHq0I+FIKbWAFvA1911JHesO35fAuu48y1uVxvLa0CUUDVjZ8pIsA1JfcmEOqhR
hhh6Ts+wpbKra1/r27ISVUzh8V2JTFYWhKaikjhJfFvpD0tfmDPny1oXUGSd6ajc
LRWXmJ9vZglEtJjpUXY6/MwIruNgNdZVX10Vg1k2JIXWftKWKR7xynFCp7Z/8eaH
yOQou6Uij6ETAjQirYOas9+CDBvNuEFTPB6z1V9tQTr0JN87n5tpFsrzODvmhVMy
W6NNcHigM0BH4qsQfp7HhDyahCxXnp9pOBYXdWJBpAzUGn6JVL6wndPCDwmU91xU
KyNtZsYS0n5a12sEF2oM/QwByVoUiNX+h/Px5JCXt+cKmLds7suyTMzBGtcnAkYG
shcGNJQ9AEinggGWaVKPeuwr8CVJ6QMuNNF8XE18Z+KefsMwJrIhULEuu3PChYeV
734QWJ92dxk2kWU4faqHo0+wafejEhRbsRZwdGwV9NbN0uFTee8W5mimkFzWZrcq
L6YKnM24YrWgF2DCGqKj7PHgh89USRpAggywUOEr+hJlbg84UrXTzmubDROXwm3o
uq/bOAi+SpVKx3fZOx20itYE0FKvD2bY6BJvZWH1aiu56EEX/PGT3c8PfzzX9wQM
tf3a6lVpJLV25CzEs7eyx3GdLxYwPhTkwlBIYYdyzXGTDeZ55pXcYs+Zk2BxyOFC
NXWH8ml8W9CuAwP1zuwg4AoQluxVcbzVedURnJLLpvsWB3Y+7ur5zfgM7K7+vVLg
VLWgwqmVnbDvjdadWOFQS1l4Kn4w88yKbxmhwH0ti6b95pzRk9flTrpd9VnUReb+
ievUWDshSkLxeUjgE56XRbqjfP2XobWmSyuzlhBv4iLWI5lcoSNs9iYHcCiKb/iN
i87w1klaZagPngBZbv1Xr4PMzNu0PwQIxdBad9AEhTygu8Aecob53TAahUvLSzdX
Cd7ULklp0Pb8otynZZzpgzC4s8EvpIITfgpxm8zl4c1yUlEwnq88VTqxVqxPZcY2
jiYfmQBvdWslyuMLhqpDhr2G5aiHXLQ3ofbf4A38uFjn4c4VzXtATOuvwdr9izDj
H/iOAA66/RJVo63+WBUtG3c2/g8nTkxXxZfiHCXHABKs2kJmN9V/Skis1rVQUZ1N
onDNgqreA6NZujD3rj13bHc1nMJzs9W1P/qKds1I7+tGJHHOoujNrSLEo1HsxzBI
Ixc+UBVBtQWzqGIZjpr7msK8q8bQte34jh4jrOnX3172f4cHjXA6jHoKigJnXVVp
rzgy9BtqJeCId2UTUeS9EPH1HTbhBzWgG8YT7FBMQT+tOrtN1/oPuczNyHDaos8/
jYh/n/136GFlw4QhwryDg/ITsbukbLjOnjEHtsfk3y0=
`pragma protect end_protected
