// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:50 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
T2sti/Tq6r3RyG1ao2fELOuwRBJYj/RxBoa1TFaQ+2BOl7P3WuYm8vLrfydaRtRa
4M1Wg14n+Haut+ZwQtz7c53SzHTc2kP4GpC67pbgi3c6C6iUFpvw0GXyvMRgBguA
sxAT1zJRcxpnYohJ4dp48FbLSJyZ6H12nfd6otaS720=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11136)
3nRw0J8qKCKMbUoxYJFW+zlxQ4UZouQhs2B9BqZzeK4cDsUHYlWYMW304hYVhXDT
2XVCh1mNtRNuPvOZvYXSKEQxC5aJVzX+nek0CGLpu0PdKdOrA6pR3y0RvqJVZFay
QU1w/nd9V7aN4lEfGjUSeArGJSL+7CK3WfkoUxMygLSZk5zoym6T7Lh+He62bZbm
GPzvvq99Oes1mNsDoyF7/AftUZeUk94rKwVi3lu1Gpg4ABH3Ys7mUw9LAtZuQkka
AX8nuC+fwz1lOKrJc792/Iy350VjIeT4Y5B5V8WOmXxmU56Tu6LHuIgeDqSmfkDt
BKRwv+a7lVFZtXoViAIjpaYK17CbIvCcv7wTikQy/xWAzoeRftjH3hT6lh2Br1MY
mPn2ZMfy3M7swCWME3YJTEm0UrJ38A0z6gWBvhFtI5omeEmSjmsx/hm3YGO3dNfG
daqzVw/ZmqK2XULGWOd+C80mf1kp+j8J0fS9wJ+hM32ne4Cts3ei1arxEbXGL0RA
bxgi9XJQgY+4/9rn/aRp8SEdTlTkG135D+t6xOZeQwkm5/XsNCvhVJH9Il/fvdFd
gcF76ZoAIzgH0RSzZ9H5eyqpoKc+avFapqJiCiavFVJJC3KcUpzz9rq1MmjoX216
a+r1DKBUNI2PvU1K/WaQERT2HM7VsbJ8k/3F6DUBhXMpr8vBX8b6fejymoA/atbc
jaYxbAR4qJ0MvqLG7i/8xuW0iud4TiFcCmH11G9BfiHCyaftxLIg12AdgJgV+4NE
f/J2IWwnAWjPaQfFTnvytMwdnS1oZR+kXNxvLiHjiswtJwyZ5SVaJ0RSBK0Nua56
EagUbmZ5fR4pJt4jbOUpF7tACX6oCJheA67eltEhOl0OS9bR+Z586IQ+6Tk/23vn
r+P4DbIeksVD/0pCnd9Ggr8Pa9zZYbabomUvntJE9GxWTD6XlVJcrWlO65lyzos8
t9Wmz8hCLDAX25WyIj6XFv/2H1c9N8cRUpx0+uIE4nxpwiN8UXnNBMwdtwQwJNvZ
YV8nFcj2thc6tnCOmx0nU7mBWHZCWI/GRPXZtQBewCVKgzPlBuH67Yqr3G6a0a9B
4RXiOCOKNQ7l+aXi112EJ99kAetX/xrJq4IWB+2fu8NAypcX12F5HFIoWHfnxoRO
p6hRonlmMJtQLNF8qE00dTU8J6DxbanVFk+xRKj4erDBkJi9wcDU6/+sTS0GaWCp
0rIsTw6P4c6iVSEYOL6f1kBpN77gB/J/E1IFaEtc0hX3Ss7z7WShoZqD+j/07T7a
81e7tRbcCeoDHDUJuK4TUR3jFqRloJVDjXqQzLJULPdcDOFsl97HAWRv3aaOn/iz
g+Zi850H8xg3Jwc/JyLWvb2gp+KYhfoMUCa72EMVP5m5Ac+wNiiKH7nWbN23Ewc1
UHTJbNJCIG0KA0OOCNmMUL3dhawjlGuH2W/lsWAhjoZyRs2KGQrHeRpUnX+Ppg3r
avTdS3cp2PSeuPh9js5nBeBozI3hwbCtuEuMKjF3qeKIWTrrOeiLJqDDQPRXb5Xn
PoJsBokzKdK2SQLwJD+SdfRkQqriICRpXbkJpy1GgMHAPJiRr4u0aZVGDhKQuqz5
iDphUFDwcZVgI5rK/4cX5LUTjPfPIh9ZGI4YoLCGWHUH8fNaMr1D1I9sgaOCfobe
lxEQxFtFk0MhS3yukuqwN7GdH0bX/00p8Gz16YLhrfCEtIzrQ3dZhFLL1N/VSkLv
ihFgRjHltDcwXd9ANHzC5gyCQqGzmWNIKrMeTQ2Nce31+C5TN7QnbkxN1X8Aijty
8Fa407pbfs28CoWytXJD0+QvO97siJqeXcpBa25p9iD7LjNh2+9hLx8j9RmJJ6t9
VfzMvbzAzj1eJC3rOmMHLFgjIkcSFbHIWaO805xUgnfaCLPilPWIXQhQd/HfMTmW
10aw/8ICOp8CX73Eo93PNjpX6J1lt0h6nWc10fUfzgu/OF+RXyb+smQTwoJzUTdZ
6YaD09Y5z4AE7p+f9GUqBaUe8J2ApcT5BjlJXccm7pXucQyAXzK7qZui/Jpam9pw
t33VJl+gDadHE2jKMDG78OIM6vTUMibx4byCpmKZtQOmab3Dx4jADWQUz5ToMPMx
/FllXUyN44D1qWltxucYSntrbnHvuzLmnMNKHshkRDl1eClg07pWVTCsmBNnuzAi
LAi7L7PSbrlDkFsBr2ef0UsjdZ8eI6/QWJce0+gwkp9N1a3ZStkudqdrnALTEb7V
k2V2D5UFXG082diCbKp+AsUVS29lQXf1mvfAPaHQYhNAi00M4H6bnaTv7iBvus3l
n9XyyUTr61eUuQW6ESl1rHrbwcoXism+Ra5bRxM0ddVOIsMnkWQibbm6KlILpTi3
K8/fy8B8DFBFqe2E9yBaXXUCUaLIAqxZ7MQjN5Ch0yjnjwGHe0vvnsAfMyRPVYrP
/loEy+xjVOqaNwR/XSQF05BUtuQ7FRzwEFa0rEVvrqd4O3Ab/BEvU4LlMFnrn4wf
I8E41jf6m7VJYcxeJCujD4pF+brgf2P6Nk/dDqQkFSMhZ2C64SMg4q45w/9D/EJq
c2oY9TXjSFz/VsqYPuZrdxKB9FPDNbo24HC5R9NHR5ImJ8Xq4mR2GhY2PoY/g7Gd
4Ub7buTJt2v8sJ0ft/oVgN4fUdYz5j9gEWG+I1SNdZaehwxh6p5W3h1ehwmRr5xG
PNmh9RBS6c0UxYFjbC/5j6Q0TzocDnqfHicSzDjmYWObAeDsGFqC2+1eikJCmlDz
OQm/gTBEwR1L4ljhO8jKx+4D0lROG31g1C+bvXh4Wy7qeMzLOVvQRwWNzne8A5Hq
lNb6G2CMRRl5epZQ9rbZFI+IXy3v1RARypGtgMG+jFy06soK8sCSKUgBDlPWH4QW
/w1sFgjlPI5TzzuRuBzS9lFoSpbuGtKLdPmBKtMsbIi4o3bBBJGuiiubCgMPjX7E
1s/i9eCw73iuW4QdNzKiUIgreFhS0c24JyQiUqBVs3QnRe+Hqp/8yEaVSyeA88wV
vBgQ1Tv4+Ec1RiJoGNvfuZetb1guY0Sa2WWAlkksnmP1cD1D5Ce0uNtTFLn1ii+2
rv99et+takPf9PSFQH3qa35rVYVvB1ar2/tKLm0zKFBP2So1rke75BMKoj7tFJ33
QYPjMOVFRNxjLh3DpybVPPQnr2LQnmCYcdnDcxTkLH5Ax34zf3HlBz5310J6COJ2
3EKmmx8Gur5W62OLC1dzZ65Mjj/8GHdTHy2+qKjLNTdt232MXboDHpz0KyyWq2x1
PoizytwQZ0+hGZhnmm5fhTl7OwNbJSy/+naTRJf2rppwcA9aBBTAhD9+NM8jORKb
UO7zg8MqYIem4p9yHIa/TwbaiAhmI5lGyuNEc4P6pEt/Q+YSrQZ9zQO/yy28BW1h
Y9Hy3ph4oEIS4EIFX1utCSRQuPKoOJ8dKwuaNF8f7cqcvUPv7jlGRQSlvRKgaBDM
e14R81te60xX5g6Ms0BznNWJ9iuDKzfeIquEnew5cG030KYfFqPGJxgnMYU7j3NN
QAZfRtM+N5sXxszNCZPWvGv5xqLMPnYGF+xkrtru5j8dVpudFFpHW5SqaXS+yi1z
Vcsoo9cJEQBm9EGBEYKnOMTv27Mrm/r5mlQeABVt65I6CQJmOUEwIKm4+CIyS0+Z
rGeVPyTssSdgsHOezfWtAVKWjS5NKpSoepRojbYtj1YdnNZgZA6kc3Rl6as+iDEX
OH3rlDtxEiU/1Tei0f1CVBavcv/Ln4/HABWxfWsSgqgXVYyIRJ09ZVx6ARQC4xkn
/v4oo8vnIZWCF0kXXWnPGJe4nP8oQtCrrIY8DTTMggivnzrmFFNg+4OJksoMl4cC
HduINutJEnTlnwMeoWV4nDm8rbMmqyxnYrPh42BoCpHBc9GKlrYNzD/6YKPA9Ga+
8czMQIPEw3zU+ykT34qWG0BBleJVcoVyQKipjrYk/Wwd6mkxRM7JNyIEb9FcJVMT
zi00SdtgZ+sIhrL5rYqx5J1MiUzI2MU48cqvYV2Bf0pPDwLI17PftKD2tUDiboME
lwZq8b9CSm1piT+BztJzISJjSvl0kIwcLCITl7bcPjmnCfn8HZA3K6U/TKozqrgH
SF9D2JCJJzByBRiq9szWbgI2bYsnxfr9OGzSR0D0Fq1sMlAXvc8iKvUUcfVbRYSd
kWRh/91neQWQHxw8ucVZfM5bOYgLb0KMMIW5HSX/kG8AzIyPqUQ7VrXehET5+Ts5
DLkSMrSggRVoqQCt3AUneAdgRaG9q12Locau5rMQldkC1n4ATz+jSYjdebJ/xGpn
SAttrom3imnF04pcWFRMzN4qlnr+yQI1aJsHry56bmgVrMVqHLwvo28OnjnT9Iw7
lSPriPo87tiutwePg/NcTbNnC7FxVeLbh3KE3pdnGBNElPFNg0JOmpS0TOXTiqFe
FN8ejmzajlvML3T793HgwEgricBQMVsVHuRkGHJG7jviO6j8vYovhpMwJWKj8lLb
Su8w3HtoMkfU5uJaXDp6i2k+aEXKdWZ+zIMSo3T2d1cTYcQSLvVKw+8MnahxXISl
88a/7LK2/goydrHzsicmHJPPQ/HB5dK34I3NT1NcY0z2AK/DQBYBjrFg/6QfK+TL
5YOlllrxGNtx3cenZXusEBBvtii2qBIEa1NQfvibYPtwdIEAoAaE28TGU1jAqfKf
IW/UA0mmHmuiPzASp9JOJbk9k1E0qXTJaOGaZQB/3IWOzJaAjK9CAqImt7TkwYQT
5VgFQmRqsNmkKYIDiRvKqN0jMXuOp08DSSyMqNq8aRYuVZ/6CzIPDfgbbL8lad8j
FiWILX0S0/z+KH6JMQ7H9pkPate1RqufeC/ueRU5V42fAT7O2IjETIjyiVhAoivV
Wu23QQeZIbnkORsauiK4rl1uO3fkVXKgT1jdrdoj0MwOxJz/2UNyohmmM3qIJfq9
LpXfj0olpQgvnJqeFoER/6UvT1zHE71EE9YsEsx32/3m0kYLJCkxArUDG0XCK3U8
eWQvgrG6k5k/OpUTcvNBmwjQCEz6LcqDL17g9QzLAGR8MzyTFBja/R41VzLw5+9S
fmVP+iKM/4HLzbXjPBgqHIFG40vvTBRuHtHZ0sbec+SYvx6X8RFCltrYjww/7kby
a6iB/7uyuOLMzpFcu0TfX8ugXx3hmACbKdmk1QDiQWQziEKlnXgsNnta95+ajDNE
WG+hlxFWpViDe4NHxgbPJBzMIRpyjTg9WgLmjPf7bgSWaiskeZV91lgE/M0R0aLW
GLJFSK0XzyCWt8tmXsY6imtDGzjRqMEgCQm8UsmOHxZbW/cGLYiQD0+faMJ7IIS5
+bdbqFanZIZzn5AyBO+mj6aYyRZDDekxpF+SuuHrOgnqnKSAuIxgM28pGWWOVJAw
GTvwXJRDzSjaHoy6YPGuOErieje6IkMYK4a+K2XjNUhQnRKuGA/9Y0H67RVN5R8T
OER3Cec9WlidMeSHPVKtyR2s7Cz+s8tnG4W+spf2lEqehqO7T+dnhY+snoarTEfv
81LOFDf3AmPxWmoSuquH4FBdo86+rMiAFRqvncHloNThybhPVnM/ZfThby7a4X9t
/LV54hilD0rWL71ZjaogKJiGxb/yj1NDDj0KC7dZKu7gsYiDiQ4z/y9BMy1U5weo
8/XyEI49Mr9HdzqrnTGi6MdIts4TCh2pse/iO/nqHEkTFNQ9MElPu0GhuPdfrQO7
iM2viGhoaz6i4kTFXIpQlQDH+fKSkU6M8Jvu/LbiA7CCvgxMA1t9qFCuRFEHJiuQ
fRVg/ZNuLU2eO78cbUCH8QXNVvQwzINFgMbR77vMukTtBHikJYyw4RYHvfOpSTkx
C8P2qr3/1NyaUJWotmpL9uXB6JgQEunKO5gfWn0w/9I6pRJ66NXt3es56N469cmk
GAp9JabLHJFrLisDwJVgK5oe4liUIgOA1lpCV8uzEYdbdVaqRk6sRRlc6zkaUzgi
IMSPS0nSqJH+oftyWQMDBB7xcTSUkqlY6TekuOlTxccsE7OzXbUQkGSgbjSUCOws
2kWPWdIwZ24IdulCTgcUCriytivUCOPCGj6+VWefAQB2uNva9NAGjaxcUvZdPIEu
9I0pMOSvSUSpDDhZg1bV46CTU4t0A1lwijnHX7WYDDsgeb8Hvf4e0eQue6hzh28V
3OECuLIij+ePSexVqjOSjjmQQ15AeDlQ0wR28XbLGfFUsRCvR8bz2+doo+X+d+oE
DIGy854Ty45GT9uhrDO6Dq++uyz/8TsqZzhWHPuzLYOx0NeXeknfMoATiv+36yaL
pRQs/5xFDNLbWszIz9TBrNu8J34KYxr1c+FR9E6L+08aAzlQfvOh+PWmZK5TfE+5
HR+Sm1QhYM0CEmRCHQUiQugUZSKv20wK8NPTlfb9fLqLV+e/IMdZHk9k0EjZUhRP
j7llHCZoub9LqPIPfdwVNzJl9OGWKt+vT7Ym/LuqE9rj2dy3UzprBE3bh6CUL/84
VShuyZCNpkKzFxv949LmWwQ8xdjAlMA/XcOu4T61xVjNjqOUN4pRYYnT6luxZGcg
qXKpPhf96ZCb2ao0mwvpCEjQujfdcEgMQr68lX5H9a7/doxuExS7+jQt35dKWErm
FvBvwi8s6mRl0cnbF7S3bvUl2vfysHaAPVAWI8PpyNgg7ijiU//94YzObFy2J2F7
6t3qRTHsDZA+Okaf6/vBcEYN0kmiGaWRpagtCjN+RzmtVeF4HFbBB8Wau59oW7UV
peZg43kg68krPrUCLisBzLfnFRKVBW44nyMYoiatcz/0Jqz7oVTxjlluDgf0SaaW
/xZ4IUZgpbuwjn9BCrwDCQlfWXArXr/mQaHHro5N4SsN7UR+VDrtilmLk3iI723K
K1NrmWs/naxf13Lrs9tpy6Dr+8FHzIxbLbq0zkvDxCWOI/EUqywCho37yMhpvbN5
frzQA2DXob1VEH4pAVr6Aqd/0o20Ah/T+n0GWc0uqhQGUksfHEz1RiObsJSLTDdX
GLUrcrx1i3Eg2OZap5wi/a4C7uUWaeS7Uzpfgc0lAC9uELa2KEt1w7xUoSNxJoxE
xvBfbaavvuvBQmQ/Ht/AsPjWSriIeIwayyzGaVQFOrJt6KnuWeDmxoQRiS7z2BaS
1sC/mKrwgLxCz4tIL5eAfetYMi8lQUK5Mzm7tA3ISJL0/WHGn8j0yPidEsDdg/gu
Z+HQ5kLQmJ/lNYhPsHa4nINVMVDqyBfFhY1+7pE3Xowt57bKpIIo5nsEmMNxBwoQ
2boy5TSfZwqkQSJVCMCeEF196cvxsv38RVXx8TRaQECWd7p2j6JsfIx8Dg3Pkw57
xa0u8+Q8PEEYE7GKE8UaC3Dvku97DqEkK8fUvOAc5oYlWmrgJTN9vg7EDY6hvu7y
JSFRyXibi6HcPLC6uf5v79Rw6kXs/1nH6S+EgeplNQKFFuW62Xtmzsy8Mz92E0v8
2EDWt96vsnj9CkPk+kL2/usp238S7wrQWWe1O3DWgXeTXLY8myixZCDEaokRD5DR
vcNX7/LGgiN6M5bGV+9ja+xY6SC33p8IqaSchPZfZ0VHB7MCXYzfy2mhsvPvhpXo
Auo+uDF1vJQNv+tSy9oyo5fJbBbilkqAf9m62Mvqcf1Q9vPiM3hcloO/e9y3ADvG
wZKYh5DinCTGORX1vke6xmqI8plvGePUHpeHywTDqqHVZ2PnHx2a2I3Tl8CABRHz
qtUVz6BRxgioAADF1yLIECte6XJstde5h+/PyJ0C3jWAEyXf7ii8E8VtpgWVdk9p
8EF1647JboRxkrCvc7ZF0o9KZixxcvEb9+/cyosiXXNIMFlbfJ7dwN3Rf4uyLPZY
QS7ZpOWcujBUneSyPyT8o8gLWQRiAXTu6Awn8Rh5Guo6N3Gec6rBgAScxHc8FnX1
qe4xLNThxUD9Yz6QZGCpqKVV2ixx9pX/ujZef+t54DhuWMW7E+ObUbUCfd/6B8qi
ysj0gh3wA6EkBmIHUc3Jedv3PZTUoSaMCKd+ZJKzxzJzqf1o9dk2bDDbwNpZUan1
7cFR0DdvcyYeA/nLUlU7huWxDS2opX4B+mVH8ysTzoUaryw56GPr2iLOkHIzH9Rz
kUw8du+Vu8eYupKIHlnclniHkPyaC+/xoQl1yjalM9kWz+SOeZGO+afmkF7+zSpx
mH7isQ24DaonQTTXsKWGAtsVwr0U8qe7kcokSYMiomf5uVHS42KJs/tzcJiZFW10
QAtHhw8AdtkZgeNZBhE1te6XJlGspJGqNZ7ZDDbmd64KlXdAxomB3e6V3wEog06C
dE4OeKBSov4PY3VGf9fxrFKkamOO6Y6+LLcY1VjsLoStaUyzn+iLQOjOR7aqY525
HXP/aAhPWV77wRnFudl1p4tJ4B9D84GS/e/R+owX1TWDnLKc1dYFicT+T0npPQ65
Uy1V0feT4B+ujH3V9eOjiJYzH/6npkCH0y8HsZYaBKl3mRzkaCc22jrDrFltLuFd
VWHRZC3eEm3cSbE5ohja+LvMEtImwjT7kliGQ/kdBbCGe7JmbjtCnSVeWg9KnGbj
WmXfCK08jUFbsr345ZRgZ0yAJJks6RN/Xp2gGKtsNG8PzF1HywVFai/+uHctIzmP
m+dzPNwYGen25Pf9rW6pDuPhRrvt+6x/2CYMcPO2SvUp1lmO3SUjU1jv88lXGYtf
I7pzrX3qEDajqmPxfKv1L3z3HGKt0geDfIokQYpcj//9kIcBXanmpjkXEqkJPuyU
gL9F5gDIWc3Zl1eqx+arymL8rCpFfSCfilVdd7R2s8zchyaNsFvB3Gwi8Z8Zh/0b
CKrrSi8tGKGuuF19uJZAjFzQyfSa3+2oBIvHfRTDXrzNrap9vUmxBtI8OUDbZyxB
IrnJLPxklmTQEVgjDCvpJXrTdSRpBPzwvI/WsuFV7NtAy55ZE0KRYGYelIUMWHEk
srX8z2NZ4hAmGVmLE6TaWvU5GLKrs0l8vuFVVKR46PmiAkVQ6ZmXy4dmI3qIjEGc
fHKS61hz/mW5xP3CJJsqGC2G47mB7GLwhaxgTzmv8x+sB59lr9Wa6glnNZqPp28z
1VNWMPVLUrAq1FmGwu7JAXcIOOqAo4vE1GNOZ1io+eDfa/20Js6fIjSqsFLyYSxR
6zyGD1hCpiF9cNMWSyBQYeXBEpmt/Vo7Kvf+Py7BI/53LDKsPbbx/qjv4EemOhn1
2TGgD0KBGeV9HmgZU3OTkixIyyby9mWEDf3yN6K2ya08OIt1FideoqdDE8IlR/jp
ZnOdQuDC4xn3/aa1e/WoEXQoYefVtwibRSKbjM4N/qnIz0jBRld4blMIKraWqaWo
IWixAsXHpHCH/5V8LzV/2EUb5z303IIcdHKeB1bkd7s+uYMmYp9HTXimySjMmO4f
pqEtFEam0viTSJ/S0qKdoxq4tUEiRcxy0oDoCH6yZOn7TC5l8yP5iAZpWSFt4+b6
fAsyDw31L4RlqdihLtLqyVvI0mCoyeD3EIJtrMlXeq0zJTyTOI13s+FQ9VU7cG27
2J6fFL4jQFrDMNMjPG0lr/yLm2esbnEDzkOeB4R52OvfHdJx6cuuY44In2Ai1T12
flbEqEQbbDCsabHp8LGLZypY9ca7frPPKTRg8SruSONJAR6nmXKakZZ1lsaoOAmz
yMX0kKIW7DHZys+MDuLPHNZBGaLyvXJN+aWfJk24+W6jH7CBwSXSBdcf5o8RQGXf
1/L6jWiOGZaF8aMmWcCDaTv+oTT5KVapOWUO3tWhrY00VSP3CeRf2AEy3O/w9QAc
svHa/l+3+xhPxDDZyoi0W74LHlV8BuxNSYZwqilF6uW2M06jrXInvZBwUKxJPgIX
ylB+g9i/P6+2KHKxhb4ghIFivxCxGFSjs6z0dwanq9IX0Vwu1et+gIYGILfigS/7
nlPndyJ206fMK/vgxSot8zzPoxPcVjg+U9WzldxFP7Geqo0EvZrDTYq9j/swWkQ+
/NeHUsl6RSQEEkxALJVnWHWbTRyUVWXLgydwM6O6jpSltRbIUmr+NSazVP+771IU
wVodFvtKJXcHQpLXl5JABQWQ+SjDHEGtaiSXP4xW2u5LiHubqpuxkonwlG0kfzJe
RP87w1FxEsSL1wwkJVFE9T8JEyRHxm0qCHLUK46j9IPlPArDzhbqVZDKJdJZ80Dd
KUVYdFKLPrpt/YRDMcCyB/SKYhQBygHioWEepVIs0GrwbgO2Di4+j5jMlIiyHgok
ZDbYbn8B2Eb7Q0+h4x1QNXGPxPTDzVSDiOSxMReUiZRiq2DyX+APsL9YbonJ+0tG
R/BULKMBkXDFNJMV2Bk3O8aWM2CFeespYwiGR8skhS1hPfDAyTcq2K96vpPwZcO6
tX83j68HC+vBFwJHa/T3b9lMbshexaG1tTHV1eZNJPy6cgjwcuk1QZUGxELwu4Np
qZ9/SWUWYmFgwwgN9nTkEml2K1JtvYZsGANzJIYU0bp+lz0nmVprdpsckg98Em/V
K/hXKy89ZF/Oo77eJqaMKJdrd6kcNihzz5cH5aq0PuGfPgqqL8I15diBmQeEEkr8
ZgMy69RkMZ5QjPu11fKZ9pXeht3hppZ73JY+kLzwY1E/jCcE1eCwa77bR7E8xB0g
Wjw6GfJ7zTOjz94NbRUzNvup/gwW5jj5M8QLunHUkTlz8xP1rfrOJZjzmEmtaFYI
rbyVFJzUF25EfvL13VvUxDgwpVD9j06xNFFyyiFkCEpAPUW5MwptCNkCYGwWbGZq
0U7TfmYUBqIA0DPH9b1j6mZfv0GVrf4QKNs6urwAjSyGmxPQJlBzG0cuELN6x5w6
gnQBodMLum28xEj4fdAeFumuJr/ZS1F+NkdfwBmovu9xmzYId4k0n6F/sVKjJ0I0
Zv5Ixk4oTgaHy9CFtQHJ97kNxzyNdZO4c6zqBdc7FSAOqj8ELam9yl65rfZskGvr
VsiNl3FT6EOqqGk0iDr0lqbOW/5qjacvdKYqX+megFa9kvkRryWDEuW9spJSiwOI
FfP71tHxaxOX3TvvGUy0/0WgzAsecxdKVOvNZ4cGDsDEND2J5L0wadHmTnjMb8yq
S7o3sp4hYqbSN4eggUT0K1FLrYl0VSPhmgHaiG26XaJJq27EZa7lT7eI3xNb4K3O
bXBveDHZmS3iPj3sEk+KOmUTEHp9sYIIoLm+KBxCwHQYtgfw7Q82vSk1EZ3lEsNm
as3vDN0ExJWXzPquL5tMUAXqyGI2lXo+cXFeAO+5NPIuS/PnlpiHvmRndzVaMs1b
eAhTnP6HyaciCRc/10km73VWSNsbgl14aNTLdKlQakMAUKRKD8kpLMgy5FX1gFPr
AZjOUAGcXjEWynabBnrW1TaSosFFJbPHskTsRtYSSyVBLiBTPfxUDh2HX48851Hk
ZnyM/sz2XAvVNzYNLPbNM2aN1Of7TxczH5oZyzBYLFmoM21hD803MC9somdPuDWA
QnXmcZg2dQ4Uzv2aolsjN3LL61+SpA1xgfZ/Wr2dD+NkUUPhFPCWVlPvGVBZmMWN
mc9ulYlxN9aVnTQHbrUXg+j4LUM2BU1VGilmk6evMbvgDgGjkOJil/B2D1dVHJNe
yhypDeWbN+aMgKFkkFu0t2RTvXg/FoxW15Kn9H7SeynAXcmQV7FqfIqWwXhAUer1
3rJzuyW1Dz4SgmKG9MrJ/gNyRhRPmuWr39Y6l3mWNysqrV4oFFYJKYob2kzGx2bk
1i//YrpXuu1QRprIqhJwvbeQN1jVL/Dvez0J3ClNwfbvkRuuZEUAErgpw0Hi6rAI
H6Px1t3lnQ4W7dPHnOrzX/Hv6+QXg0/qSnr6zuBrdVNQhJcNSzdzX/D48lLhKZIP
+AJMASTA6viEsx5RdnBzITuFAu3c5mOjkNfyBzFY5GTtBjlV2Xt6Qdve3hXeP/sk
avPEwACHwJleB/JIH5YJbHZab9xULPqXru/5RC8z5JSjZfYsXlF36hcPlrAknLx9
F6TbkXe7jQYiUC6/rgNaxCHpxC6Ay9QwC0PnOyrbva1P2IZcakh6RH+pTgo+EXft
+jOPFDj7MrU4wbgaHcxh/MxdcFGTbNEy7glr7rQu3g4uXILngMhx0IOKltabM1Mc
8I6l7iJYezSINCYJag5YM8IZYSSstDpEjXLukn1B/FP9Lxn+5fGtrDBbu2BLEclN
faW4WATk3L0cMtntX1JSZ1R1kLc5Skm2TMS2HUf8WBczNE5hAZxeZsZVa0bywD5p
GacQts4rswChXa5l/s2yu1gaAD2JadJuoBujXn7TalAy8CoMXXh9ek6N260jTST4
6phXn45yKYSJrrTQx5TyortZ37iol9R3tUT2GagsWsAZ78LrvpuP1AvlWPF2U/gE
RgxdXbQQhhSTJXxnBJ3/jXjgmpp7c9NfJvOygiSduU+fMm2/ypn1npEkSTyUfj3b
nYMpzCyoUzlV9qXU3IVe3dXu3LFW+lTks6tTtYq0EtZoX5oFgKNTV+rruDoj5VTu
pHlWwlXdHNcA2B+PF63nQXJkDk2qar0CIsbgqwtT+gdyloHEv7siRD5TX25aiZxh
9JbuAUyuhNybozZyG8o3fYMTuX1ysiC2QTDRR1zoRklRY+rdfQOFFTGfx/PLIJPv
FGpi/E4L1maE8t8gk0d/KDOVa8qLvpvlj1lZXvuPLB5lRuHlVn/PEngNVFvsl1Ge
RrnLS5CBM1OB8jxYdfB/+1dJFGCPQT3z+fd+TTk3EzWK6bC1NsBcIjwXmv3hCjnX
i4NJtIo1iIcQW/02Bgp7onRCzSskUA4gq1vKLSS/b6Pw//pXdtSpsuRG0U/LDqVk
NXInkJA41mI5gCkQv33NURFSrWlDtsff2jpex7ZZjcCUM0uZ8yyUEzdnmIShJ94Y
Lyb/YhC1JCNkaHzIDRvbzzHbIKnOH3AAj2nDjOyHS9A0wZAKW8NVCiYLh92J2raw
kNtDGCJca9cmoICn+aumwCcZ8zI4kpKzcIBB24Qt/RcXKZB/7gyB0rJP9sYZQkt7
LtIAmErczJntNZNcPQtjsfGl8wDCyk+yU5mGRZl9LU5se4OL5klLHErCXOYiRkV6
mnhTELGu7kadt6uLT/NrACprQh9IY5yD+YRCFvAQy3QWJ4vd+Ict/7Cbh2oEt1NZ
WM6/xjnsE52XwMpMYxbtEBNFdeDxR7qBXdznfnXG5J+jAm+cyomNwxJtzGIvrqVU
YbBBOO1pUhLMGLqoLFv4mGPAWNzc+LD+e2zf+fB0XQJQnSHBopOEOtnymXqJQTe5
1XaqbjIsll4lZIosQbbqcX0zg/fZlasvc2cNE//EYcE/1DxbepEu/IdMOju8jeI6
PiXEMWsE7qkGjpAghnKMireyG8U4MBh944OvypEmbJwNiKpFfBFM/korSe01XLNL
p+Fgu6k6iXRIc5Qe9HG1zy6uAg96bRVWEcxQomqGcBtZVYsj90fnfs8Vo4sxtBpA
IkDtamRDBxDg1ZDhcN6m1Vf/eBnC4Rj/RGKNdZn9MzwL7DvbPCUQiaggBGKGLr7y
7Tmxellpr6ih4o3CH2Omek4SVYZGC9EnznUaiOO4sXttUIb/PbWUuXBq147U5e9T
IlpiBEO3J7h+AgyULiTz6v116lKdABj0OyKVZQMzEAwdCX+m9Sq7HTp0Thn+xas3
ouhO+ZV7D+XIK3pUqU1SumlrTplEQn5iSNyiXsZeJ7CrjiU5Ghlwa+EwJ+80SYmE
oevTlq/sJXAQt9c9MesxWMiaeFG63R4Itx5iyLQ38auC9PatCwqVGomsB6mL1Akx
XnHVDeTVxqN6F588R9+Jg5tH8GE8NaxedsJLYheWz32fbr50unr8xzLikHj6j+/y
KJB2PLJD36FJlQTfX7MhcIcSQioDiUWQtr0WEH9LkKU7cfW/7TawTo/w5EO8BNDI
NLt697rCtf/RDkZ8eOng0qDy/Gi0mDZqmcZm3cbKVeFKZtjkzIh2CWOmYIZGweYw
Nz0flpPBMYpSNdyXWeAPRcUyONRLUNvXB6cVk0bFnsF5s7wUqMD9y9kE3Owq5FAM
EadtoPaQPXXV50P/wgi5ERySo+aOfNGqAK5MeNi0C+WwtiSA65LarxadMzQm+DQP
6zYBdYHlQAINdETg+ilLJbmHVOeQpk0FDyKIoCSEiJhdc3P7wtFbPzeMV4EvXco1
htMEFuavCi4PN1aOMBQlF2apZjosNMNC1CuM4H8M4h4r6Qvoy5/H4TF1uK8F6YoY
j/i3Ozd5bVimhW02i4LvUou3S/XlesnhK8mLwmB6vodA1cKE4fbr07K21JKXh13Y
p1r4l0xq136+ZmrVQLmR1V7UYp53wA6OFpSAiE3SLfCfE4UlEZLZWxq9V+y6pBeW
gA1YFbefL/MQb7Rr+BzeQ3qOQRwrqRQchNRBGVS20nrVEVof6gTt37pSbU6ZQX8W
om7dLYwjcSDtySixUXlBqi2OYOWMTN3wvYrx0CQUASSdWcpLN4itfdidh/7UfwYi
PunveBKPV5TMc0CtozV6gQ8a70LRe82kuSWm+WZHhzL0TbEFcbYVDMruRNbshRW/
vj4Dra/kYygtXQTZXliMoJP/UyAtT9HnP+6Gjaz8BFWQ5tAFkW99PtBWJBBi6ckI
vR6w6Og0AiaIKZU848m7NlXJvK3tAs0ilFeQ1+ehhuBnIvz9rasE2PqOAndKopj3
OVZJxnJovhpRKwq7O4akCtmFOb56yS9MOFvoDaWRa0qjFJQ9d/P6ftEnGaC3oVi8
I+XWGi9WVPq3agJcbD8A6UlaC67LHwZEABt/yOmcfE+/4/7Rpa9RF88odqr8uF/T
A5zpNyHpP0R6wf0w8wOG+yb0oUa9a1edbnAYODHyyFDjm1bE2H67NPoPIrUGPIMX
Excn4h0T5kTuDbnqNLRrSBS4xXyQK/nHjxe67etF2x8xAQKs5Aw6a3k/sBUUaC+e
`pragma protect end_protected
