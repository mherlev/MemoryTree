// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
`pragma protect begin_protected
`pragma protect author="Altera"
`pragma protect key_keyowner="VCS"
`pragma protect key_keyname="VCS001"
`pragma protect key_method="VCS003"
`pragma protect encoding=(enctype="uuencode",bytes=200         )
`pragma protect key_block
H?Z#(IP(8 1*":4)2?XVVA(/^0/SMKK!X!\I4_'FAU@)N$$2?^-AAF@  
H:,>?9+@<21<C-ASN[&5B1JU[=,FQ_FF-CE[J( 4:$6#RBN6,?)_+OP  
H8'C#9AP8GR=K,8DCB&Y\-F=BZ:-/*>Z5;\#4E(S"L+^8VX@=,7I9FP  
HH@[078&.[G#5"S?-XP?*K;(PRKJ,#L$<KB!4R+R4"?'6VMCN8BFS1   
H,?HH=HNK:-UGJJ6W3'8ST(5@(TWTJK!9BWTVLDGZ7V<Z'QJD+OD4%   
`pragma protect encoding=(enctype="uuencode",bytes=13744       )
`pragma protect data_method="aes128-cbc"
`pragma protect data_block
@AU$IX:1E.\)?4%NJ)'=X%G AWB@7RK,2@[$WRF[9!W\ 
@]T/1@!Y$-BB*V\NA<!AZ@2 KI#FNV4$<XF7\/T<-(2, 
@& !3 I_.L@P831G1>-^B<C\]$3<.3IS6&L?/8B63UJ0 
@#,H._1=60_-$""M &2;51I4W5W@*"<<:-V/<SZ-*2-H 
@RS?38MQT+DX)E"K1-6C9CGVDJ=#SMS,16"(%F!%EXO@ 
@2L"P]6._&EU<AQ_#2C1DT!:$S0SQK3]<1088 ;'U4 T 
@\!U:UEY"T0+$B?R/F/'G-/?Z6]W@:3*B[VSE(%8!NGH 
@ Q(+7T(#2D^(N4;'S\K2UX8B;_0/I!&Q3O,N:JKGE<8 
@_?9/R9.X=-\-L6KVW5?XVY5&EC.C0:%8!U#ZI[P>.)H 
@GC^< E.^#^BUMI]BZ+BT>I(3R<FLXE1)4.D,J(I6M   
@A-KV_&+4W#[31YFPFH^HR4\[B%RS0>3I^X,VF5E>!D0 
@_\"\J!) *-GMOS N1EK*DCC4^UM5='8.JN KZ9=&23P 
@AR:DR9_N#-59%GKNT',]^;\=!< Y2Y=(@@X9.$AI)8< 
@1!YQI! D]&2!7E+7ZDPJV!,+3MB#QV/FU!Q6/VL_!30 
@E.Z0$OM_:VG$2[3KI8)EF9SS:X^:YFZ%")W,30"KXZ  
@5XK&YR.$]V L]IUF_=Y\FJ!H29U^HN)1V 13XP3@?H$ 
@E_^T2[EN&FQ,W7IN7.!=7F*?T/6%*UHX2L^HRZ8E=$  
@RK>4?B=%5-G5-&<F&6FZU8<;@-W%=&4 "?%RW.)"<0L 
@#Q0?Z6#/IH^=5CO+IT6B^:]5Q(7AQ%?_]',40Q:;E:P 
@/1,.#K*,$)$VLCG'B5/5XWZ8"X\%>(](F./^*LD(P.T 
@ M)LHK&T-:CQB6A.LW<&#BTE%[8-B,<A<E4A*_=OY5( 
@ J59N=BV%ZC)L,SV6056</F8%ZPQMP7_73PLJ,)BH,T 
@J8D\*W060.(E;(1_;+O2E-$Q/5".+!8/$(,]YP1%?C\ 
@MV/0?_C>\E0>65]8!KX[-VAJ2?!MZ..66*!7[L)_+*  
@K2]EBTS'U>B'^$V59N,4.>P7E-XW.T=F^]T.4%4#Y.  
@^FNW=L8#9I,SXLO);&03F;/='[6>(YV]" S+()F.!<P 
@-,PP^U:BEZ3:-<* D4\!<X/!DO??>WL9D6?H0I4BL"X 
@S#JH/O?N*GE0)@.2:"E2> 8$3J1&;.FN*1F_NWF0I6  
@9%$KQQ_IG"^Z^PTC]XN;6Z=GE1_F^6;\JBGZ$Q,CZ)0 
@4\GQ5J'\[E0*GZ'G>\H,)JJEB?)]) %9'$P%^U71DUX 
@,^^=I!D_%C^J_J>S^!"L&K+HRQ5WZP7X0/<]D@\3= H 
@T&'YFBZOQ90IR'%6.U(I";U9?9 %Z:%R!>(#G6@SLJ  
@FVN9QU-P>A318U[D![2Y56DD4$<N)7CH%<RI8CCN&U( 
@;"F87R':__2(\3 B,?;DN6ZIX-/(=9*/,(&XIM:G]KL 
@G(1&TW;BZC8%PD$'66-DAQ $6*,8A>/;:W',ZK1SLXH 
@7=3@K,(NO3O#]8.'?5$?I31%^57V S91.%=,[PAY?T( 
@H!=[ "2VH-VLD1*W/XG_KU$)W=I9:G]">K >.V4?]C0 
@HL1UBM+4]QL"@427K=JQ2AXH'8D9<W"6,',;)W$T@9T 
@2I<=>; P).FS+@I!&HE+[/M^KNK'"&UX*NWS8M/UNGT 
@5'YWK2K"_F_Q!3\-XGR;HM?$>>TO$/[.[6E\(9#?^8( 
@YNOE:-3VSJ[D;-CZY$HDZF7OAN@V=0%K4<PBQ35\*U( 
@JA'PR/KXV=U0K8&WO\:(.B-,%L1'6!DJ"O<P7E8TLIT 
@S?#+*JQ]'0PGI-C0=618"V<--?"VD_<E;WFI7!O56%< 
@%?P'6)P1?URANEEUL$X9,=+LS]W2G##<[-C.2E'0"ZL 
@H$ L:8MV+#'X'OHH@^*-$[/@\*J(Q!XY29GLYU-NB($ 
@0KN6J3)E+.L1RMZB'HY9;0)MFFD.L37R<%J1(K"W?^( 
@>XBWF(>:J 71DSB.RL(UA:JV:&X[;=%JX/F;G6W.:$D 
@;G>+*GSO!OI@0SZ(>*CK## A/G[LY[MC;O%TZ76=;KX 
@O_71*5O:K'$/[*2&PP[7=XELBENI;!I;<C9H<X_2_F< 
@QL)E)$-Y;]XD3#8M7$=V,S34*J,/.J]])4"["Z85/+X 
@E'33Q=#=R)VR3'ZT*,R8RBV(98=82(/?K:*YV Q0P#H 
@?+AM=CM0;=EB0D*_[^-2NU$!RP4#Z%D0/$\HWZ(K,=0 
@.IPH0EAW"6G=@!!V!.X!-$8LW$J5]G4Z!#MAER*2M7  
@KVR3 7)[(<F.R/2>48N>R!FU,CW )PX$XB<T6$UY=<P 
@_-1)@7>5<?'M FX0\ &0G&$G9F7.$0B^P$/HN_R3"'0 
@6"4>9SV"W<QY ;$M7UVGO:_.O*C*_M2T);QVHS>$>5, 
@+:MT-:D0_JMM?8-J^P[6:FOQ!F>O3)D[4@R]\^]WW?, 
@:QRKGG6G/:YJ? !$WBAK%-RBF*\ K#W3!0<)T!+(524 
@OB2OZ1;;(EL$QM?>6XW*$Y@]2U/OPA27_<EQ/UG 0I$ 
@7=8S%\S=GGMWM0^.!)^<0,NQ0P;S]SYQ&4,;UY/!Y%D 
@>8K1Y#[.S$ OT_6RS<OL3H<2Y*ZHHXCJX"HS&(2@<'T 
@]^QO&]J411K#8%9G1^#?80S#9+O>@[2I%WK=;*B]?/8 
@D8XLD'X"QX3RQ!+/+;L$=TVPU/@6D5OQT%JKZB5B!T$ 
@W3UZBL43K:3+G .#BM'W*I08^\F0F30]H'\_<A+]6(X 
@3%W#+;]B4L25)X2^<@&OP@[N'OZ.E;W[YG("H<?US[0 
@V,F[1B4XUKJF-0%P,W" BA'SW#35M&JTM8<<\51E+?@ 
@.CCN(:Q]2ES8=<N2OW,4C#EXYZL<W+$/BI.JMVQS!TT 
@0(MA2 \V@-$E#Y1Y;EZ? \A=8B:.&20^>2Y9A6O.(B8 
@<N0EH!FIX+3$J37!H+DK-A0$,U=R#\AAD--5-('.BK< 
@_<+"R=F7<P0?O2#%BTP@*!JH%;(W=H'W;K<@+XVC;&( 
@/5'%90Z[I&Y^Z,[6_(HN,\?$BA*PZO":-X#V!CQZTW4 
@^<&>&<"*0T&'K7?'A?T<8W]UR.)H+J\FM:L940ARI[< 
@TQ02^Y OI_Z8:HN3U>EES!Q"Y4BF\5#;]5:(6E8YA2( 
@ZFL<79Z85-31"(GD!4"*[JS%E6(4<W[C"/<-JW?M*DD 
@ -%DEV_;'U%P#5AL^+*'0 [%]1CON:R@^F8JU!WN0N4 
@@/1_W<ZD?UI_$;V8O*8?N38*S6!".J_@_&L4@CNU!M0 
@A/JF<X4JUKY 2-J?OX)$;DEVJT@F,?T#X,?Y#,DY<Y4 
@#6-T04266T.'0'MF6Y^16U&123:!VPTYJC'QA#TW^!< 
@AR@A[?N_&#I-\F]Q!"YJ.2#7.&YV\VB\M9WY;@M8L2P 
@,UD"G65N.5&K?F4'Y3@YKG9RK@2ZD!(5&J_Q>A#/EL8 
@_KJ&321QJ,W^C'%/F8",PBO?+C/B&VF1,XT#@3SJ.GH 
@0A?RM\R@^QE:@+WM''<(6RHZ>!8ZF*:W2>(D:/@#W]X 
@NU)4/X/;-&S3)?*P@AMH*^WTN^82MX0>D;]2 RW7 ]8 
@4Q9QU*3^#=8 "E+A+0B)GF&_S66&CU^X'?DVVXY,(U0 
@8JUF:+-,4*V*Z]!LD;6@?2C^JSJ?O3'S /TP1$X+&CT 
@'FYXC938 +71R?G7C6E">+@XY&/.T*U#(XQ?LY1#HA@ 
@AZ?%1GM7L8B;_IS-*IJHZ'FL,+'O!Z!PMMJ7=0/6Y_P 
@)K<:@:=&MFY&3W%<M;+@["^!&*%MN:28XUX"^3+:C[X 
@+FGIL @P?2^#ZFF"+R/O,)%;A0PN%]9LXN\Z04R4[C$ 
@<N0'I/&%<-99W?LW0+YA 0P%_%S;1-WWM9T$2E#?*MX 
@6#+)H++JWR+E)[Q:FS-F@KMN2SHW2Z.?L4R\BW$&P_8 
@.$(]Z:(BI+D6;<@K&(4D 4[ZEDS '!J.\P&FL]83P<D 
@7QOLX8'S&NKJ4O 2PP6/=F4KQ#A=#&2X#3G*=M*% ;@ 
@X&?H4N:0 /%+O29^U3N];J>:!=.-S2!8;3&BY]_I+Y@ 
@QJ=2.H($SYVS1E^9WTZ)EI]<\>L , 9C*GX% ,DZ5$( 
@JS_MTX23Y U@#6XL,-SU#WT&>?5[GXK]KT1N6BZI)'4 
@F33$F:TC05@]EHLGL_EL]G-CZ@3R'X4'Q)@!P7<,1KH 
@@* 44MXKB;YOO*]YQ&96/*G*V-=#5N\\%QRLUF.EQLP 
@3]*T*M+@)&8[MKZ([NO*NS+@H@1+ ;X ;;&JH%WM;)L 
@3^D5C&OI00[DW_7M*QX@A/K=)P\]IA/O2./6*N+\/!4 
@5[1BBD5O"V?"7"M:4XC&:(#KZ8!O%13%RK4Y$PR6T*X 
@<L5KLF]@U0^AC)>R>/21+C+7TZ3V+F?*<F'Y.<DO! @ 
@[31WO%.?E7,C@N/#W:<%*Y'C^4,E$Z\4[6+BG_3_>8  
@FS\N_3UNUF8:L2!J?$FJE;'XA/3]$PJD,GC59B*+*U( 
@B3C5#=$?<?O5X8 J2=Q!XW]@[MFCUAQ(0!Z.<[D_X@  
@4#503@\%8.S*U]^R$@%?LYNBX'G3*;?J),^^PX:C^RP 
@12;<QP=Y(*C-OKS9QK?G1$8<RM%Z4V;K4#>@)78Q#_( 
@H%"@@@(\O,.Q8*UK@^)CO0I?6:D!::&,D 0-D-7.?_P 
@5IQ7S)?0U5!.M2O5Y@3HL_Z),;/UAW/.AWWT5U=KV^D 
@29]5-;("M0+*T*S+:,YFO/60F?6%-N@&0]C!Y@1<U;L 
@C/=8PHBQ G[*JXSG2?QH0,_!V>.B]"RZE.R2^&H,-'$ 
@Y(RSHO;OD[:4]GKS/_"B(5HRG4!B#12*( 8\%.Y[XDX 
@')TOC7L9O?_28O*GY%X"1$I/"4)T?P[6 #EIM5P-IS, 
@8$^EPO2S<CR%"/G)6Y7LF+UR,EO#BJ;$;B10-5I;BS  
@I::MVI9>QM!.ADJE6DA-^KL&(RVU.IAJYV-X[QUXN3D 
@8=8#8R)#>^KRP$UIR)PU,50X >]NERR[5B,%C[-I_PX 
@V0?DC-BV/G1.+-!H1Y*E"O$X8E+U!4/;S'QO.^7Q?O( 
@6IMV"(;N!W5\Y^=8W25<)8"$CZ\P06V6$&P^:Y.A)9\ 
@NK&4#??Z>=; &<4U0,I]6M4"((,@#%YC0'C;*&XHZQ$ 
@[2VGWTEY"-[N_:(JK:W+*342]:6]#5YY+IS&(54#'%L 
@)Z#VBH <[,P *B(B/*-)S8/23' >:BNAXY*)QV*GV'( 
@*%[4Y.P<NO_8$!D9O+S%H^J%9:B9C6F^Q5:,?N$/%:, 
@;)12&?976[F\38@=S7O0!8=#X43/F)(7C)GH[A0%^(X 
@(U)0#.C8&9JX\ZCO(&#-_2"ROH7KCX- J'<'1^NUTY$ 
@MI%7=Q&S4]"DMC"N4:; ?'-2I\N)4.[X1:2:[/X[B'D 
@9\/F<\I!(P9+B-:0F&(0(_GUE1I$TC]#Y!ZL4AE7VMH 
@G4LAZ#O_EV^62KRCJ ,B9#ZOJ[ S3?:&Y03!('K.4%( 
@/CPS3T?JIYU0>"O]1TGK&^?MM)B_Y+F(I9@Z>W>G(EH 
@%W1=V.I0@3ZR)^<SQ'GQ0O-GHDI7%L'7"L^E$<C<T)D 
@\?7U;F941$C"FB_R5+P_21IUDY#GAEMYTC^6.UX$ @P 
@EQX8M\ 1O.TY A!\I:N$CF+)LN4_A]\.H[I@RDH]"6P 
@D9%O\V.Y8CTX(B+FV\$)0,CJ(E(!4<^C5X@EEE:KBHP 
@D4-XO6CHN:WH(7>9&PH/(0G&)#:BZ3" KY35AXA:RO4 
@V1A-@;&6<-=&*.'[I!>=/;3F]:LV712KPN)V)."?L_< 
@!947<Z(#Y@K''4/O<:K^:7% /:_!< ":AZEYO,!]+?T 
@X-@\#S"HRZ=)DS8(9NSN1Z],\?&,<AG:\0-&*KT,UIL 
@EU\[N6RDH\K$A< S^<>HKS[[+>&&.E&D,;T2KI)NEY4 
@?X 619W$M'C1J]3O26XPG;#]JYNOY(']!^0[LFS\)9  
@D:) ^6=DVH$J%/+&>*16EC7_IG%!QKOE#S@H\L:!AV  
@Y57*C*ZB]E(1:["=R)V*U.\!^?4,N@".0Q6V5M0//+0 
@;T-ZH.,TTF,#Y 96@<$>@@YC8.A5//G]>7_N7=^=U/$ 
@D)ZI3,I26?^C]=B@*-50'K=M,TF [Y):; P[8N%OE_8 
@4#W"U6$X<3UDY#$TF9],4WFUIG6@PBJ];G5A[B"Z.S  
@9X/P2(D.Y MO6^8_DZXTG?%L$H;'8.IR/\&Z6"8-(E@ 
@[2U%-K% ;UE!6&R?5B@;\[:MG?;O8FWVJ].^V0XIYQ4 
@BJ4B!<2 'W&D]/KS@ O)1,C)^S@ 4K>7I),,DO%WP"D 
@<"0A#0GN[A@-]*Z7/!KFTDR1\]M2H")QD YB0T$4C!  
@W9TNS@50QSI\1 'X=H$8.AU@[TZ/Y^TNYWD!SG&G/IT 
@"#(R=(UK)"CB'X:7V=USA!'WXM9,'U;3FVP65SH:MG( 
@X(JG<%M^<!RYD/.HI]V:])_>%F(P&,Z2!P6Z->Z(?S  
@H(3)S[E;Z;EQ)*%+(>V?^1&LQS3" %JU+#YRZ);!O%\ 
@R)GS^6T'-"&PTWWPI9P&/R-&NC/M(J2;C@E=&>5ZGS, 
@N;XO2@/4Y'M<RYX0/T\Y&F'G:N@TB#4&]H#Z(2U4#04 
@DR$M]N&X W@7=4F ?-TU QXYJDMRD5%;B,2AJ(C2?P8 
@)U%C7&/BHDK\_V%<V7=+_^U'6!:7HIXQ#;D3XS.*?HT 
@*TV-R\Y:/9[ Q_ 0#'F+3U3*DJVN]&$9P2-@W!\+M$T 
@M3$"S0QKN(/@1.6T]0.QD_(X8^/;W:/-I"N$K2O&P 8 
@M#%Z78ETSP@RNDR&55T<@X)WDK)E,>5&<V8/WW&]0>( 
@H8NA!JW\_E.Z%C.2\W*/9I<!)0A(P(#CT>BB,.O,:'T 
@ T9MH,[>12Q/%:)"K<6"H;!9U>07%;U;79H.RT]F" 0 
@X%QC4=#Z,0DD8_$[0+HP#!\-\S42@ Y7HT2Z.EJAIS8 
@$C4CFK&=1N)^AN%W!5YDO_SGJ"[1045=8XYT"QW.\T\ 
@5YBVX)F4! 2!N?Q/6;;S&Z;P'F"<\W3820>(7.T&_$0 
@>*70S41A)G:724\"C'H.S>I%B[QFM-XHE8C]HD]V=)( 
@:O:QUQNLIY6W ]%7Y\=FV]L%]=B2K+TV:ES.CT[A.50 
@-S8 621R +F']GEB5"G@@&LL4#%?3QZY!+)])+L%'TX 
@OZ]#P_NOW!;Q_Z'HM#6P:P<W":9US/^BUAZ?C4>"H;( 
@#\N0TDD(VA%;#ULHM(E;@;: W$D-B_7,HTG\@S"Q<&\ 
@;AEC5!N2KZ -%*FS=LZ!T-9$_@G3!]<R&OU,QW&YR$4 
@;DF$+V'5 ;T5O<88,U#(<975BD)44C^RI54FI'MP@2  
@P[*\JU4^#O!UL'Z'?8]KI.?2=SE-\XSU'W()]LO'7RL 
@%,R)01$Q^VIT"]B)4(N#SS%V]'3[C(!4!/T$7X8K&F, 
@O6SV*:PLEL"$ 0%.S>Y0*7?'!VZL<NO.>,1 V&45SX< 
@,_9OT87[8#VH/KE@T%+RD3#?_NTDT>G805>!EY!2 GH 
@YS!4Q<+LCNR2A37D)EQE=H-0W[01?)SYA&<8]#75,Q@ 
@TG4YU6/Q&QU+K= _[S34(=LJ,,'L#HHLA+/2J"\CR]4 
@P!DA,S<)0[#OH;^0)B[,.#=7]R?Z**2/8X>L'US^L#$ 
@!0)LP9*R1!'O]<:IM(G!,)Z/&[L=_-RT*AP*^BB+_F, 
@&OIO'V*S-_.$POVI-V$/O<7X VO\&:VRNN2F>N?RU:, 
@]PRO*Q6]"3_X8]%$0!G,TF8RBY5;;O0 X*#2\V7L*A\ 
@DQ[ZR)F(Q$9=(>L+%-HW]T,%T-/Q 1=V#B=_?P]T!8L 
@5>_0> [HG[%YLIU[OL3U=K=N,<'!R 94(>N1_ZI A?L 
@FA<X[A)VAD&V<SROUS*#VJ8F^X.U,9L?07&?S6YAB"$ 
@[A+'J^\H%G6N9@)OT.8MVP:9M)_>Q]:]W1<LKT0UT8L 
@/,4I#BS#Z_YFR^1DVC.Y>_\](2<&%W!HCX/P]10IX$H 
@-Y=6T3JQ0YB6C$5E,2:)$J?W6S4U/E <5J,T)7T<"I< 
@3D(CI[) 9SPSS.]L"SMZLKIM,S;?T.KF(XY@PQV1,14 
@]B_EVAG^UUA,]:='?.->5DU8HYNG\9V98H?=B;;#V5( 
@\X+(],W$*J3F9'9S).1QA'UR4-5VF5C3CTND/W5$T$, 
@]L\&+<1\W)(5^!U"JTVBK;\QN\215M*,K=:M0(\#+8P 
@<TI=S\6$"TL/AZKX1^LD ZAL"6@=E($O,K>Y3T<6P)X 
@D@[T.N52[@2^:5_0OAT.7SED"X(%^;>PS%4GRY05L\T 
@F-L1:Y('E]2(M^SN&QW2+3-O5-#U0*AE$[?[>[RW_10 
@(\S^%72-2,Y"*'P*MD'ES9W*U SA%I1_ &7X9->P"]H 
@%8!E5G-NVR_G*S#&3RW1 J:>6[>?.=17^CA;7<0PGSD 
@'0]:9<'=/^@9*3\;]HRJC'-)K.P3_X=_9,9DN.YC<>, 
@N'XI2J!+C?FKZD:#:-6JBKF+VN+6FM^^NB;3"R"TO"D 
@4G"/.?_R-!-A7%SE'Y;V3GCEXFH>5Y*7'(<K*&.K8OD 
@&( >=\ IM^\_JQ850S3W2L#?S[B1%,"Z#GQ:MK@8P'D 
@1]R#/]PT3T-P3HP=$;\%;A2'TSF,;&>G[N'J@S<.FRD 
@0UXC.&" LUT8BB//)5YMIUR3>#X=;+.@-5PIPY/..*@ 
@7'LDX7E+PQVZ] Y<*ZUXT]F?V)XK N.SQ %"$!/:W%L 
@7[XI!N:[ ?D3*]K5ZROH$=15LU@,K'P$*JFJTH.F+SX 
@M^Z6L<4VW#D9EH>(>U7!0HGF\'E,Y=N@,SG/N0*D%KP 
@-XHI%B4)UP9)A>]=M\_ S/ */7D,VK N>R=4'#3(L'$ 
@;E)*=K'5GY:H%3)VBA3#$:$/;MX9,GGN)THPP+\>Q,L 
@]EI_IWYU"2ZP<17Z7+:KN,+5%NZ8#EK3A8\O=U+AW#H 
@W^(#5]6-D"FT>LG9C=!L([962<K9Q<9TCFQ<J8A[ER0 
@49$=2"@4\%IT((CNTM 2-7-*X'@:.MJ,Y&K;-HJF"^$ 
@<O4,4^-.@0)\^$H25<:$;$U))_2J",(_#D(ET>#S?,D 
@7&!K:75:<.*1E!L5:S6 QZ2'><SA$A EPH,].CQ FB< 
@Q1YQ6 *'3^7'(@$M-\CU*AER)V.'#LIOFHQ&,XHQ1], 
@$5PS5_8J/LP7WZ>JP3A3:\B7O_]9&2==$!NI:JOCX<< 
@.3R"]7LJ$QL ?U(X0LGSPL4X"\ .E85DUY6XG(/&+>D 
@FMU6,Q(82(1Z[ZG;+J*;6.+!E]$%X(X&)^S_#/B\O0D 
@:7S;1&VYA4,$])[01<\Q1#>FZL19B<:O.+(_< M;:E( 
@XXZAT?>O80T'!3^T:?A[YA>W_=+.A[\M;!CV= #$I:$ 
@9D,Z04J\,5I%%0(7\%@$!\+"EXFN&U4MP@X-G>_ZW!D 
@-:$81KCPF/QHG0A+N&,7PTIZ865\>\?#+9"WTM+RF_X 
@J(N]2T^KGI;[$TUTOW([5NBO[4(JZ%07YDV%4*=002L 
@1/P*FZ&,""W..6+==% E,! DY2M@->=T!<6(&A[-PN, 
@_-3<W4:8LE'QO"F^<L%GRZ+!:7CHEBX5/D6T R;8C,L 
@.9X-T/3/P<XW68RYN4,GA30"T!]^[SKME3?"^B!8M^L 
@U\6"-6=_)'/:]6:%9-8\M1>52!6')45XXUJMKVNKQU4 
@<+4) 5I&I17YTT8WS2Q5,:S"X!#$JICO ?6:GK//8)4 
@/T*#SBVS '7*MLZA976?(.\M]V%=M=+2F%4-J\-5)/L 
@K'#-IZH+HO>OK3B.GV+YQDV9Q/?H:[6XS&L:)JIX)?P 
@A'EW2A*U-,IH&=!O$_N7BR9W'PUW?AQQ<5B8GC322V( 
@+H_+K@NH:")9<1<3-1B#D?QCY]LX,O#S(RZ]Y-FB=2$ 
@=2?"%YC(P*B#S/5=BAB1!0ALOIT%AS0YROF8)C/YH)0 
@\%>^WGW$P=.,(H57VK8'NKA*-M(S?2VQ+UQ^JB'&N>\ 
@WDE!EP/LYIVAMI3(&P[<W$)W_O0=3'* T((^F6=!]M  
@XPO*?5!R>#EZ8OX-FC;DK$]A+N"_@$J^T]09&J0DLAX 
@.BA"9&;'EIS!]M#5)];8UJB6RDPGLA,K1#*;)SZ=MND 
@I:WBS+N@1/5:^;50O:J)*"9W%0]0,L?.>0\$K^,RD+( 
@F7'=FB'"[<)XLWA+DO8R=+85?94AH8)<5E0)^S(*@<< 
@-?7\K3YYQ); .KPOE]?OKP@,@;<8 V[4/\'D6@<-2AT 
@XD#L_.1"4 =L5U(1QGRE$:P"V!^EWPBV*7,V*IS36^  
@0Z0J?_\<XUSX.Y:'% ^OF+ ^3CM_$L2$^(*_WZA%W5X 
@S/&!! ?*?!S_'QP;4UMC4 3N!WH+<8GQ-#ZCQBGL^W$ 
@SX>&40;C4#^1=.5C<X/-#6U'NQU@<MLXIT\@L>RBGN\ 
@->X2J"SZU^!++:M*EHGV*9.9&HG:88F/G1,"35US+54 
@N'&N!T#"6<\-8O6KQ:3'L5.>?/*$E5IG_ZA+_NIN>>L 
@,Q][5S:8N97)KL4RIT,H*SSH-AY596_--1WHR*>>M*, 
@L?-6$Y;\#W ,J@5W<**A*?M=KJ<RFR7<F6Q<3A_92M4 
@V-K;.)M&TWO^43T8"^[$6 &3 C1:2B[T,X>)&?8R"HL 
@.8&Z_5JXQV'])).PKV7:$/=HL(GN;'"H_,NJ)$^&VMD 
@4HJ;O(9-<*2&YAWZ%]TUND9@"*=I.XI@F/5.#!((ENX 
@.;V&O=[ <K-6F*[*F'S50%2V6 EQ%W, G=X8+'N#N'\ 
@@>;@9/$,B!F#E"Y%-U<6WE5=WEN\$NGG=&V$(*7QZOD 
@2:MHH]A"-Q]@I#<R(N@>1.+)1?*ULL+;,&?.9JW"L9H 
@@#^U_ULY;CRES:7T:,1X44D@U1K)<*8]3K7U@9)_PP8 
@'<V@[8XVNY6#6_\XVQ[P(+Z+8NG9$ML0V0?P9F3494L 
@?#H#,I4/XIR.W54R?[_"/SAU;V@V,84=7]KL+;0'K(@ 
@U5Y@KAY+*GPYO 5V#2R<"0]7<0_=[ZV]35(J7=/SC,( 
@_@Q9T*-OF?*2[L,TN9-NA_Z*^C(4\>30#V>LJ05%O%, 
@."1K0U"Z0_4^;6$#(S,4E#8*+!"!V%:.>&9?JM023/  
@\?;S:I[Y"-X"!^9^.JFOC*T;PJK!Y.49M82 7A))"$D 
@:#M;]CO?>>9P;:R3ILT[]+7,3(\<1T[S<B(#CP44[=H 
@ 8. DK%/8Z?-J(*8\.G0'$+-+_H&IZY_I,K\3-;G!T< 
@'*_\QEZAJ#E)'XW!>O%7SK>/*O[FR%.7]0WC1+J'F+D 
@R[3%QKHUQ:'\C>]3S*(033>#S#=B<C><.EO6[RLED3, 
@YTB;O$0-VE"$UU>/? S"D3M$XEZ1,D:8O"-(&I>]*8L 
@O!67<))103_K3NH9F;A&L1D>/%=NL#N3D?_*[NI]IN  
@2PG,W?W*+?Y#:M?<^YT@@V0MA_>#9?J"D9!VV?C_)K  
@Q4PO91]F>@Q*#LB@SX[<E'3L91KBOSDDN&#HS_!HU/P 
@>2FU-E$_JA?:__G:1'$=:'DVIC2L9MOY_W2G&FD?H;L 
@B%"#,<S6LUNVQ,BWI $J9U$CC=AQP?8ZXZVY[MK+R<H 
@(@N#X0M*$DX<*,])S1<0QL+CHU[%P# -GC5_DL9+D_P 
@$MYN=<N](S()*$O$DI'8,L?*,8QL0>,/*29!9ND5F;4 
@D][RT4D-S,1<T6#^T*RX!OO5/(VV;CG/0[J:+4[CR[( 
@'__A&N@.M]R5L8!5?*R-F O4<DG9'T_OBR_24H<JF!@ 
@TBYZVO(E1]_@54JWH7_C-B6=+VAX^&3WRBVZ$\5<F!@ 
@UF98L;D;&G!E%NZ&B.7O7*IQI1;D.MYM<@P.LYM)V"D 
@'515[Q67./7#<PC@,)FYU7&)4C]E4PFBH2BFH5A$I T 
@;:]]S#>+:0KE6TW2.93"E0@^&X1OFG/93>T6*>+=M@8 
@8-$?84PEDL,Y+_3Z54)DOI:%H+2)? S,(&B/>T+89,, 
@>EH@+@_A'&HP4?K[)4518"#)?@D.:+IA)JL3&ZK/C4< 
@;-;U:A+=6=29QS_Y/6I%330;O$."+7GX*K1N&!.R87( 
@K7)M788LEQ[\]8*XBU#G<=;DX%>%'Q%B'D5_=TX <I$ 
@\/^T.9 1+SJ_NO>E9L;BN9MI6;$I02\C6Y%"D%%L\W< 
@C5!S[ <**=#]AI-1/"_!%1#:?#W4E/5_28@+?Q1M-$( 
@W5NU_,T W/<YVZ7,/BF@::M7FR#\-2>7-<E]IC:X=0< 
@3($T_OR4WC_TWE^.>H(,>F\_H4I;2BH.;JN%'38_.1$ 
@7N$UF*R%YH8>5492)Y'YSOJSL2V=4HK_^8_B8V%.:"4 
@9R B2E_6W?ST<;?O7DV34--;)7EW=";<G>1^6H*J>=\ 
@K^'*>H #%Q4-C1A.FF)?(-C5Z!%M$WMKEKV<"1A:_*H 
@&\%D7$E[;G2)>=2G+I/8;FHAC:\CMTA'*LM?<3[[6=T 
@)-T'4 R[ >\"_G3T=\"'<M".]Q>L%40\$W%2^)<\@,T 
@G;L':[D#D]'LC:*-"0:-GQ^7#=',314XQ"FJ*V[3GXL 
@3\^Q()N:D?]<7:^8#YO!8WM*F8TL$@XA?##9P4%M:+T 
@?N@69F\QC!X<+D79+XX66 A8M?DW,)(1-.GF;/8YB&X 
@K>G%U#G-LWK(49M]J*V&$T<!&<Y1M\1AN5R$F^^3QA, 
@!MZ/ U+@:Y"I;-V=$'AO02>(.H/9C5SCL$KO;<[Q\@, 
@X_[H\ AS;X?V>6R*O$V2[712K[&_\5+OBE3>WD9G1P@ 
@-V+Q<P2]O5:795(RM: 56&? %BS1-KGN5K6%D(F%KJT 
@O[0RN&",TD^35Y9GUUQ+$I4!$\[($Z'<(1;,9PYO(PP 
@4%9M(E3BQCP*G^_1MZADB.FG:&6N>4&-B:/?193I74$ 
@1?(J:3_8.0?K97#G:KYWHMC)%U0.:F6:M"NLWJL6<1, 
@>^#-.]R0S<YYE#DOE_"J2V>&GZI'U= \/LO7P\60!M@ 
@'+F4HWT'-*$HMWI+1L0[_#)PBB8B!;=R"TKN @6Q#DX 
@.W"^7UL&:>2A#><G-R7O!A^A()EO(.;810/<\6KBYT  
@AUH"Y@M:,.*KS6STLH31 Z98JIR9%VC.)$Q^>H;,[UD 
@_W]02C>U, ,ONR^5*J]B.RQJC'%(;.]]Y&H7_(YN60\ 
@*WX@I70&I 'UJ*>L/U99IP.]75&0T+W.@!?&Y.E82@( 
@XG9TJP_\LS.];J\Z;,A01NNY8,!X_ @MLAR85:<S$$< 
@$G-J 9.X44!$U;@VM#U/[Q<LIF%&-H]ID1K..DMS:[4 
@591:P503B9%O:$&J=:9^Y%@ZB"W2I]7?>$:LYM2;'>( 
@ N4K%Y\J<T.C>03A.?YS/7$8F:S-9R8-(6=E6T#2-Z  
@SKV-CA[KIO2VNP- )=E+=EYZ:!.YQ(TWC??H/@P!F$  
@DW$M6>^(+H! EA@YOJ&)&*<R$JHLN8S7MK+^J#G24I, 
@@KQR .=A]8F[?A5<,.7,V)EQ]7JMR@>1T?'#&H&^$%< 
@=+%;>/$UPK:.8(!9")0",;ZZE@P"[,C6FT4;BS:2EW  
@>M)W-CVW4/<-UD1*@)IHF'@AA_-XY9<"-ZC%]<"66V8 
@056\6)1"7'N5]*KP>!.RL=+H1]ZIL2_?/)0D0Z?M>TP 
@*__[,R(V@HS!_HO0;MXQ/#>X4::GHV2LN3.:#AH&BYX 
@\YFRZT2LPN(G_>OLH?$!<!P#M!A"6E7%@LL9+?[T]V0 
@9%RMT[W2;M?0/FC]M2 A/04<=Z&1FM7A2S%"97TMM X 
@ZE(5]A+W-H;MVM.N@G;ZH4R>;R4(]1EI[S7=Z,8_1<@ 
@A_965\Y)? L$TUH"K4)RB]*7""3+&:!_141(FF5P;D@ 
@3@PPK_Z1A3]49IT46V ),07;!HX(<0V=X1&$F"ENJ8\ 
@4VZHD23[6D@MS+7(5&=;NOYN.VP^=?:.K\QFMV[^W'T 
@SDN2Q:4Z30'??=)$8XH'$.>'<5^U^"5PU%_OI+1P"Y, 
@>C_3%612%W<75W31XY3CAA1&^V"T7W]0 O"!E+F-W1X 
@.LF59%*4%4+=[WQ,VIX85",M69J*\[WB<2MG^+K:JW$ 
@ *129FS&[!=>OP7)=?K!287(5*<)K%9/L\[SKUWX000 
@)(2U^&D59UEN(P"Y0%$ZHQ.)J5!]OEL*97?K,]/C^U, 
@S7,\$.?L*-N$3_%Z0B%^GJ[-V4D)4<'NR%R: V9T'ZT 
@VY!,=79X%9#"726B[^#"D*+6I?EOJ[[5J%*%'2/GX98 
@N92T#LS!B6]DI<=+70F7SP6%Z\A<1+8KTKGP"G$,0L$ 
@\-.IRO"T"49/219;OU!R+!_3EF6\JA,W T5A8!/SQ   
@JOS0YI)UUMWIONCL>O&&Q==-L$I7W]W<8OD#I+=JWU8 
@_(Y%%['^@8?_SM RR@@Y<[,?32?-5)TEE*8 YE-A(#8 
@H5L>*_OW;CP#@K'_*5%B'<XQ/^F8LWSC=UBGQB=ZB:  
@]T&[SK+#%__Z!J6"I)F5CA$? +"43>9JXK,KH-50@54 
@#2CW\E=41U[0)2LTP@@?6>-D39[".14B*B^%Q8<L16< 
@X/S?_JW1.^,^*C*4?N_LI9O_XC^>$>;;0?MJ^&+]Z-  
@BD=$HP(A),_FZV9/?%B4KYLP8V?A_DSBO]!,8;+*\24 
@U1@I?WS0=// @S5<-FUE. >XE<DSQH:.BS\[4K=(R\@ 
@#A6PT3Q0RV&-Q^3#2#(,^Z(M_P3XHDIZP"113%<T&K  
@\%+7>0343'Y=0DG?$K.M)WA^A-#U9_W)FTMQ5W[ B,  
@%N%D3RZ*J$[,,!!:5,>P&GI$8=ICNL#\$R?F7*",(80 
@LA9XV,R0D)PJCG[4:IIZ:=F9%] :()UL(UR\L;\=)UL 
@M/VO19\HW"2+%%>DD)W=E9KTZU*L:O,OTV@4;796/L0 
@%'^7JH;H"I^3B@/0\)M4"Q->*B0URPP6?,P+S8)G$I< 
@3K"MUALY+Y-Y=*K=XU7KG2%&58-V8*(<Y%.6*0NW%R( 
@ X<U*-YU8(%N_CUC;8/E?0Z)?W>"A0A9W?)ZF\LB0!X 
@@&4.PX$ZRI[2?*JFGT+XO/994K5> E)26;'YQX<_<L$ 
@$)KG#X^R%LM#UQL18-P%QP5'J]!^5Z]8$=/FG+^C(9L 
@*AJHB'1UQ=XD0TMZN2"O6'3964W5!+,T*P(T>[YGQ$0 
@T 7L\!&@<EV&K"T]K>2H12E=)FI6KEX+6$Y\[=.J1W\ 
@TQ\\*ZM5WQ/6E^]D2>^0\3XBUE35,.2ZX+=A_"J"WBD 
@:[I#8W;"-^/SE_KZ-@6JOO6JPLVL<I"#89\;?[&711  
@2(:2BXT^5UWO((@ZJ<R,(-9Y>IGXVJ<A^7Z\0(3Q,OP 
@$5VTX?D=MRKY^ -*E:7AY0[SPDA(*L+4PRZ6:RLI26P 
@!2)IAUKS[O=:XK]YVU<[C&'2)YMY&I"7$N.UH#=UW)$ 
@KRX@"B2]F/;93RDDK4[7<RI=F'GJHSL=H]YZ#LK>P9L 
@LUI#-Y@&%)PHN%%*,I8<5@P8)V50<X8C@@6^!*6RG14 
@\])[EVPV!^3>X&YB"8TT/"0ZEZ426V&S$-=W.^'JP?P 
@[  NJCC39@_4>C9I['(E5QA<C* R7QB+ J&I1)VF:6$ 
@ 54=M:AE&BTGPO6I?I'Y@^A^?BBP9DWL2[#QR>*EK0@ 
@J>;XACE$-IZ:HW86D\KI(;V,%]KGS3H--IPAK(R.2CL 
@)>/ SM\83S+DHU\V/G#<C*9/DU67L'151,H^$H)Z%*  
@?-YY7+\/;I9BOUC[K]7<_$*,S\DL#EC9$_0U<031D/  
@R-^&0*Z\&T,ZK<IUBJ:?UYMO_3$8,3'1^^9,U#5G0X@ 
@AR'OH>#9>7R0#B'^-B\&C5S2_P*HJ=:+MS(<B2/!E&@ 
@_JI5NAPC/U>D0AK64CQYV$KX),N8"MSF;O6?B*'^K?4 
@@4BPA\&'%H305@.&1_=#ON15M8Q+)2J<U59L!2(@8C@ 
@WOP/GRO3PALUORD1?SMZ23+I/:GQ$/)8AGIA86T4P#P 
@X514.66%C1[JJ9.23TM\,RL4@6]15'5M2 V9)S3]_80 
@<OK1)6TRS1RN&:2VQ4B0V<2\\#M'11+0C'O\'=,!?Q0 
@^*.K $XGUHUZ?]8G9C4B%RX%KWO@E@5V3-2QEJ_2+0H 
@U>QL\(&(_0K(I"<BFBI#:UO'_G,E#O)L,S%SM>'OC_4 
@]S679)5PT6'ZU4NW"H:$S'=Y9'/;L"RI5[X;EMUCPD( 
@2Z@O]7MK?HQTANA#ZYR*R;G _TIQI?ES,9$F\ZV-5C< 
@/K'>#4I&2AK0](>SK/[-4%0BG^XGXJA)YXY=@?/A(U\ 
@&?O+7>^VHO1FO*R@F8O8A.Y]?N$2Y$YWI2##(\EF\88 
@[G (&9+<\Z$':M\CJ;2OE%WO"-."<RK%ZQ(,5&VSC%@ 
@'TT0_74^3"1D#&N9*I-BP:V#/B9S-WG)!?1;NV)/&G$ 
@<:ME%X09V'2, ZS27F!P_>ZUU;UF!''C+EMH]UF1-PP 
@+U9W%&%*$A?1E38FKVJ!U";\NQ<, 2AOM#A5X7JY5OT 
@#L -8(2I"4"$450SX+LPBXB5,.!1/XFTC\R-YQ4J 'X 
@=53XB&)<@BCWY5#)C\UEZ[1<L1KG@-,FO^ $@=PKCW@ 
@5;6[ I_?JW>1US><8[H7^)-74'- *_>86WXVJ[W#8=, 
@0V^6?XEN":)D)(\+X(P0'UIZ+))^4UXWJ'G.YW/AY>0 
@N0VDWXHIQ:D?W6=%?_SJ^=-[0F$@SR$,[*3FNW%+AA  
@P?*%#&S<LOY\^(- 2<S#!W;3A+-10)\>-$_&K?W !5\ 
@^AQ?[2<*\0T]Y:#\TP<J[E!KKOK6<9O/&]?;[C,"'S8 
@EX .";^T1K7!JJP$T):;9KD<12.2$N1$\.^PU1 W]XT 
@1K[8@@OM^9&:5UC/279>$57XNTM::O.QM79AZ&LSWPP 
@A]P>\*RC];D&=IB_&@R0)JQUAAUZ\9PB"[I54&=DD1H 
@9.4#EDHMWVMS%F\P/'QP0-'P#$ZA,)I$*RB'@LH[J&8 
@%-=N=W )_(+O\STQ0'/"Q!?8575("LFJDMN*&< A6_T 
@(T+2H5?BHOC.P]F0,UC.LPF!XL0]DP-(%KJB+<SS@?X 
@WI=6V/[$7JDGAH_]7DKU;MW0@?VVWI1-S5(-$\;Y:/  
@V2GUS%^&J_E"&]RO@GND+IS._'LO"7$1U5Z7+%$ *"T 
@_); ;/]:YA$YE5O?[N?&O))P^4?UTU!DSNW3'7PI_DT 
@U9Z>X'BB,P'598<8PWCN3/D FYZ84_RJ7WUE0YMY@>< 
@!\Q,#)XT4%^XU\7U%^G!+>S6^S7$,G,]1<83H<[)(-T 
@%B>."05;@O.(YB]U%V"/3QTL)'L!-JY5RLBCQ"WD!"\ 
@%CQ&[^]8=PL,!4<VT@I?KHZX%'L-N;;,<C1R)W.JC@( 
@&'9K\CZ"^V+:Z7/-),^FUDH)XJ68GF32"VD<*LG]GT( 
@G6&]^T//D;$S>DC&G=%+RI_??Q_*O';AVO98#(I*<T0 
@K?VQ1M7VNL; ]C4'V^_U71A)_)]-!<S<N<_W5O!D/O< 
@I8$A<^JZ/-F!9*(#Z7V; VQ-JSQV[Z LEB2Y *80^SH 
@4GYW!VUHO$ H6]>]VJDU;)/=A[P%SV#FR7CGM BY9R  
@891V(JGQ16VGF0U^S!CHMR?:0[<[&[XM90\VI4]"0OL 
@M1YCCU$XFV:(*>C3"U+F"<1P>9WCP\&%2B 2\J?XQ%P 
@]&?5[KU9,YR*+,$6S<>PJ.]:XH;];9$Y!8>^#682Q-P 
@KC\:R&W#_EHW*25H56J]/EQA9).E8:.S1<A-Y"1^MLX 
@@W+\]T*+R^5]TCQ:O*/;[6G4P6$P&++-79S.O6Z;(.  
@*C.)H1>TC%)5H[S-"Q/8" H'!"?9=!L2FZLF))JP0V@ 
@'^,WE)+1A+'L0\\SO2B2]87Z9-/6WT7>YJZ"O31D#Y$ 
@&$OFN&"O'IOU2D#K:E /UJ606;>NNJ&&UB32=# UF$L 
@^^"X\1GOU^2F+V;V\,@G&>4A=6&C73)[C OD%83RO3  
@E"%P%<$^R4])U+)+A*_05B< ]^WZKTQS+OVL^E:_6AT 
@Y'S1A#5.)QC;TJ44'-0,TF8Z2+4__C7;BV>'5N9KU@H 
@QP!J/A"=-561ME!YJB@-$TCU*M?=-"Y\:]SLF;T,M*  
@2;;71[/?$7GV!Q5%^![:"@.4!65;>^VT>@W2IK*N/-8 
@T.,2V$]<S*P^5X[>R6.P.^9J[%4IE!R683UAM7POD9( 
@J8B>C0$APV5 "QP'<.AEZ5DL(+6]+$P.1YI538GN:"\ 
@X5!EZ&IXU!?;OJAJ@9F;X#685!=RNW*D"<G<+'27QED 
@5%K$;,L<.BJ=VO+)L4-H.&@(O7U )+_^H)-+@]PXA:8 
@]N<FDY61^80^-$L<]D$I,,MH _2<3WES0\60G?T?D*, 
@4\4@X=R*T=TJ@T/Q4 T[6?XIV>+M0 :@E*+LQ"&F[C< 
@UX!4ENXFP<"E\G;7P.,05[:>D?:<8EJ&O:BM)$L@8E  
@C5B'>Z]5\SYFCFO*7M$:&>5T;L1TB#%"[FQ$=B=YLJ, 
@5?1,B1_CS! 8PRT=%(?,-.Y[-$%#AWF@PLI7RU(@.;( 
@NIV&AF])*HE VG1>ZB-Q0EP(Z7E44F*/>363)XM+D/@ 
0I=9"P&XJVTZ:=!%->X<J30  
`pragma protect end_protected
