// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:47 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
IgRgmW4tXUI/jvWfUn6ghSdroINi2c35gOMn/2oWpJL7nJKUitE5NOd55tMz0kLl
lpeqybXTf8uwfP3Qw60agdGgn+Qr1Q3mFsYceyS0oP4DN5oQmDWWO12ThP9N6BdD
B5brj8/N4KGaQMCGpL2AyV57wFiaoVIzZtDR34H9eSM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28752)
FDAWvxJhwiSsFMbytdgZB2PrUEBeJ6FvM3N1tEJpb7q9rJruH7zQrbAD8TGXIh6W
zb8f5gTuFRmMc0dXu/yGut5Yowfjlf+PZKgL54E3sPoOPPSReDLF1JgmcryEjdvD
whERZk2p6sLxnSq+jMox/AUNEfpBUCBKvZzWvK3fvbom4NghrUvXDZ4cMNYLv1Yv
pcnfdNdgOjJaGdPSGE5gWjjln643vHXLnrrf3Vr6Z/es2+AgKjhGwMJA43qF4TSZ
63aYCPocRZXdwb9QSLlJClxxk9ImS2t8Oxw+Y98c2ltrhe8zuJhsXXe9+6GQwixB
HzfCNXF5yba166kp+fgqfRcr++ZaConvzddfbPpN2aEyQR8xcXFmdX7wTVymPOMV
Khk8C0Tp6ddgOqg3Iiiv9MKh+mvl8QQp4cwRKMWG6iB3AOmIF4t57YsJV6s7FMhm
itmebnd/DO5uaV63lPD4guQjUnQ28hClNNzW8MERuoxGyuSJNLIUyWcTDP5jqn8J
bbMJYzchONOjdFgO9D+9zzqMGLI+R6YPxIKpxM0BJTpVho2zk+BGIARm2Goo96UX
l17WQmoAjZ8Gtl0Yu/tnZaIwJJk55zfaRsLwASEyoS6XdfnQlS0oYUviqVfDQ86f
z+Yodikq1MEE9U8mRY37Moo1dQFSUZH0VjtYX1u8Y7th+edF6VDmezK8ElxS59kS
8E8FZ9ssl+4eopF1vNNFZb/PBpBFSUvfaztbIe8/Pskn9I8B8Iok/5dABTv/ilEm
akO7qeu8+z9i4cwB7Y62siw7n/NmgIteAuxjblLKZaHyd2ApeqG/UQoGN9YKUY96
sEmkfbxuko3Z4omLQopdNT1d7n35c3x1moy2OE2yx0GKWpPDdjIX+3aHzD/FaboW
Pse/eewyd+OLaTBhR+k+CtBVf7Y+OycR8PsEhCd7aZBdSq2QsM95ZcCBNWhQYFcv
+6RosDrp5UaHbuoJvN2I1d5znwYlPlkXxaDJShXAxmB1KvXPWBtq8dtQZiZXfrmh
H3x/9W1fahqMTKXpcRs5QypckZUy2/vBh+pYDUlURGyhV2DMhV1cmW74IN1dW4Ac
aZObQTRbECrn/6qMvBYDv2qE7XZMTwYRu5x/8ImFvVbacI3O5ibLCFbqNQDqK+rE
pUORS/4w74AlL0ZPlLm6+rntOxkstsDh7YHeEIQfPfvaqwV13tZ4TUK+8RIpEGvY
aR3zpTGFkPMuTtD+DQEXU+MqQyyZYJxoJJV+Vmwdhb7E0FE+I1oQGLOQnxPMdwW5
jGSEBgR2IZCoJg37Mg6/am7kmfQ52cuvtUIAEubh59GqTXA8tmgM6I3NHcSHokBI
deDmTbNJT3044AnRBwwS4wvXTKsmX9uTEhNb6rGb3We5LsQh0mc3gl+kkY0eUcG/
lV/S5Sz6PZtRB6XmNMAxJXzhFXfY6J0cl0FUz8WiNrmDM23BmI0bC2KdhTlv753e
afBtMt9S0EQ5DmXYRSNkorA/LEhdKQMVHtqpfCouyCIJDsLG91KfhFMJs27WEwqY
vri3Yjy5gwmSJVMnVOcDiUQsDMO8JXhT7is3H1Zi39krSlbX0Z1MXYwjVJE/PWyx
AMQDBFTb3cA8SwFTAMQMQt4j81Behdz5c3pFSuh5CB8PkQQWK0+b/zhQHVK4NKmZ
vMJM9k81RYvY8sOTKy7+30i4kx9ZGT+q0GrNGZaCp6w4rfhGwoKx/yFP4esUf9pX
cK1EVvnY53k/wm9To6c3DQd8EQwMJcJX2SkIFbk/zPMMQ0XOVnwyYduOUiWixigB
sbNg/Lkpg4ocwZvf8c5ifGxEQuDS0RXkfhTqXpB7MhP0GliVsUdtGdRPFj5+iclj
m3cBBxFE/8uKmhaSl39dHSLVVWJKFJYGdNmiZvWPCH0UpjwPNc/3OoQyJdFRb7EZ
R4j4OUlSg85ZB5gVY7BbzFXTC3vVsaJuNWD9Efh/NI3/yx/DG1DhcM0GSWBHsPbX
tbicxKCCPtOWTW3aq1Zh5Q77WSCr/XGAK50VecZ5PNwN9Id6X1f1ZwXn+13xjEla
Edp9is27TLPVbZNEMEYkbXsdjgr+lS8JEwUbbyO9oF3n6U4h/FnTUt5ns/MhJuhi
sNixiJktXgOdRgrQatSJ5koUyaaCHzwPM1lh2LjbICWAoAFKwiT0TRTspFqlPxz3
8kVkzC4RvO8tdKCrCqfMXWIxIigbkjTfGnk4tLzDVD9c6xDO5gCda0F1M50vOjLR
fXli0gsi2qIVBUg5nhwbgisP0IhmzFiZK94DU6U+CUAEhCKBeRISoXkyP489D15u
ZR6Am2WxFxAcvgLDljelGflAVdOgpKT4uzDbfq5NqqMxzGsl+i8TFRtgpz+i9kYE
XNqTbec6DzrYpKn1HcrPAYYPMcsBxRWcl3zzpCRVIw/Tc2E1Ge7If+hhGAhUkw+s
EoP3UGAVOqC2eJJRyEwoJQPIRPFxgP4yOnW9c+k1a/C5CoTFCseGe0+64fizVshW
f0ocXreCeROR1kIAYFgV2JjzhcB4ez8fHv52MLJxttFIenvHop2ORcXQ9foAepPf
nh4ra7/ZLq8cPWVr8S4bdLljd9Q3568zJu8RmdmBtislngCQ9HW3n7y//nIgknef
uiI86YAzU/6l+fqsElAWDLLjB1aCA3eJHzzwytfVKlnFxLXSxbOf1aZ2m0yuRsj+
faQAruktSsoM6U6NR+amYNvr7EjDBx1QGs0lXesEXRevmzhNMwBhEn0I+EtH+cTU
E5kgLpUTxzML/V9n1a6Ip8UcUkiIXOVhGJ47SfbiqDh0qp2NDr/aXPeuA4YSNi55
uXHeHd5bBKx2YhiWdOEC2Tfrl1ovGVxGqJLMZvWF659mqWx9LgU8C/mDvGIA3+5J
Deb4zg5vjpqX10SP50hjHBn11fNtFmw8/sSQYJGRdIJgv/7ASJ8jlcVgCFwKxtNp
AwYXLMnJeR0RtEgwtIX/IRzAxmwXNuvuLvLFaEzB3VVbvMVlT0p1GurMcw9dJ3HS
3RAIIhPnSOdIA7ztTt1nQXWzTyUQe2eexJ0gl+GW9uWPWr1P7DZdIMp8qr8yoQbw
fr6a+oXSxU4tpM1WwOYoMkLdyl/FeYGgTSchQuh4JTwUpoeD0BNMGS3TekriXuT/
OPVXgUr0yV4hJHgQYsO1UxhsD3WBv6qxapJtjt0IhFD2m3CzIk0L3+tAnT5oM3VM
Vq1ZFZghIcwlyt59N6DE2wF/QMFJulOrkQH1wFY+kHe6W9IKXNcYXIbo0DNHOvQr
bIkgoON6M3CGd2MwTmHRJ0yWDewEQg+HehcJ45R1s0YsiUqLDMXUpGOQ9xNOkoeF
Mm88BwY/ojh/gnuj/Y8KSNl9GyWYdQM3EnOYgjZ7g1d/gfGvnoMotpkuYsCNFfSF
7lmwiy4nTqu7bkm3R8PcGJ7kut3THJvRkSw6DPaxSoOS7zHbL7w7K61cebiAHSiI
H+3QtNs0OJ6Z/PCtY/B1s+dKJJWrUT9fM+1bMxfwgcBKxUINNqSQrhxQbh41Gn0x
UKyBZ8v3kMs+iJOaJZxRPvGabpAMbtisbdySkwmBwlHbx4wYEAeAsf9U2E/ZDAvM
5ngHeU8HMgeGSQML72iJ0J0o8kBi2ITM8+PSDgOSeX814LdQIhVJXQ6Xh/WLxjpp
j0BVC3dRMQr67FVFuziRrMJ5+nuQP0F7qCUvNq8VGEZ7wD8yiYhnycfYURZWJo4B
dJ8qDQkXreQ2f72WUOZ6Kjr+kbII+iQshelBL3dX82S8b5yoJ8KDT4jtH4mPAmVc
MlQNeI1HjVaAEq6Nj/XQUqxdrN8cztmL2JHzE7zNYFlWaqwpf3kspzLwnX8GepNo
1dFDgtx/0HJDoR7kybumSSi/wIpCvQMk0Aqx2zXleUMHDS83Mq0SXPZ7b5OYrVWv
829cwxR1IQTSGcLrutanMiNCIxbIlTax0p/iotjZJVXYxe53veW8FjBBsOUaht42
/Uq05weAgKh0ioFccaruxBfszeMmf/aR3Nx4iUxhX1XJrVXFfiCnbZUbmr/QbHod
mFyHYP6T05hpsFN+h/WThPjwkY14GcanfOswj2v7i8mjrPACvGxvRk8m+KR887hV
3XEdYpQQ/7LyUnmzf5dDvNY6kzF9nXyNnhhDlezQmubz/ASk+JHGe7VyzqAC8VdO
autRvdBmuxiHMKL4FWl1Y/Mi8HAfnZPGOdyy3NrmDgrIuOna9mWz7HtBB1UiLJ7c
2/3pKbUENMeqbjk21zqlggWCJSidC7dybpMOVa+0fX3ZlPJR3h2MbLarpsES+4Rz
fr/3UGPWuF49Y18sHIqEGgv91nhqU5xEr5I4GqlwqS2mOUN+VCtTzk8HNUmjHRZE
rpmaKlrnzR09AEJWhAuWEvxRIP/5l9mrrUjiph2ldsQXrMrWk+ju2M92IObYCaRr
xVKfTs1Lly7lYodyVdxSS0XxqqE03os9mnMDT6ri3M2XbMUs/if5wUG0GV6+TZMC
wpbXXOUAd6yQfQRiwwDEmsJpQQxYEx0GgANPuAKw9QBpPG8/3Ym5vg9iePQEQJMY
UwsC7Tf2pVHewa7FSrkkayX05IsuIFqeahYxz4cK87We6AZP2lQXCKns0v9hbf75
E1PB2iaH2EOwVnb91dg1CKDKc9q1dTYZKg9CbetGSYAOITovvND0vJIX+gaxme97
CLVrqRIgZIRS41XDcrSqEcoWmzxRiR7+K9wLBy68j3HObHFJSqHvxFvR+MQR4Eaz
qh9/IGfmOfic40naLbNsfOpW0v0nx1dQZLfFAKAQyad6U+45cnGfpuFAr/WRieSq
l+E7x6MdytlW38id/alDXxgJAtJF8sxsMpm7lie2F3I6orzzHNLR5aD2rcZ9EKQF
R5+nqfKlmoiI6v29t2/OefzdOg2Px1Q/mKLLSOe83fcy01LodPr1OI00isTxg9gp
8W7EOwL3bWhvqdm0U5vULstXhj3ysvp0EZ3Xv/lbH6f/s5cz8jXcRLaOG8K5AUIC
B2f5xac4q98nilC1enD2gHGg0x0qI2XkqduRbvJLDQZ9ZyjxshZZyNJGHFKyM/0K
obwy1nN8RwtCa4CNUcMgdd9NPpF2sJgDg8AkU0Zn5U1cMii83/8Dd2E17SEvwUSR
c9oBgss+kfY1NVSKf5PZ+mKIjBelhr8gorxTUoq8tNWIC4nkTTIQ/NxNFjnwqON6
esf0Mdjpm8A76v+f9VvuS8QlUx0t+ltQqFFUOgyeV0rIlzdsOK2lMh5XSTAb9gYp
Vpp8t3VR99EpZgFyuH2rbouYgz9AM+JmB188zSo3EN39cDQOY33voSv6drsgt47r
kdK78/pFymw6YiQfXi1Rwj2ME3A0k78NB03RYoZ4nsiWZ7Cm1Vq6CMNpyuwYk80B
oin6gHvIvmGkFlTfapF1WwtshRMBWm/OZuWTMWG8IJaxMyQznsiIBi+cTpe6C9y1
hsn60FEe6iYVeMDnc2pjCXOIEiRLeE/ha+/MuKS/wrbbGSE1gm2Jl48WpFYpQNa3
+VM8BWGU4OBTRhyM1ms1HMqszlLeZfm4JDxvT+ufcgmcnIWUTpaaAz/SA0pf27ok
nYD/i4+pdnyUyilenpqJUKe5uHS6sbd04YoiSs4lIyNJd2EItekY0CZhaK1zManc
YmQ34ElHD1rGZT2PBf2EEsHY2lZ00excUFVy0zGJZL4TW+WDrunxOg9FXvx2iuOy
R9h9pYrM0p7D9Gpu88R9uBJfgSyNQ0Ik+4zR5XWWYMMHHGENaNNNZNw8M91FyIvo
9MFv6a0YtKe1Z4wnLGfqLMHqFmbhegZ/bsRCzg+NBa5XvlT14S9/nOGyIq0XdcaJ
2q8aSw8Uyt3i27GaXzjKjM2eyAT83SzHJYC9FfivYNbV5to/gz94GjeYa8REnNTF
VksOM86PpUlYPonUTkQzQD4lzBHh8JyzWUvFjFwqS7NVquLAq52M05gDYIkLojcD
bnoVD5kto2eT5m59dAwUN4BV1i927Wz12sgY2VH7HRelTmDZ5As+moocUxS0m6zx
JPkVFc+7yT/2oJjR7xOD4V8VfwSwwwS9ijgl4KbE222nx7Kme+7aOjb/fYsKcVRc
0F7Ni2im0eXdfeqP5bosVvsWR8CsoxO9Nq6XrH5GtIYz9st0WKObqKeqd8NXpq5t
Xd2iXddnkiWQRJ+NPqv6Ej9iXQOAT9gKYdzHGU83OnEKXyENVuVJVRIcDw0wlx2A
m2LP/ivV/iDAJ7FMZF2bYmvudrGCrntEURx/TZ1OZXeeNYLhKH33dnxfCvREZyrK
Sei2syKDo+/RwJAS3csT8XkpxxdCOEKlFswZSD9w2/a/PBzywYq7coUBBhNDrCXM
QCAiZOT+nDp5d7FyAhRjDuFa3oJr6Txft+u63vwWuaGVyH2b5MpECmhfZWh/CckA
gG2NE+LISYmnteQD5XggXH2NQgCGelJa3CPoWgDJzDE2Yu9kus2NS14Bx2GIeqXD
CvGSsgtFPXr0wgiPctb2zHCOaV2uq8cl5rX76Y9KUDHasuF9Ms9J7kVr7mqfif63
ShriQdzlhIUQkHDunofRnYTppr8xvVlymAGPiPIoK/HxU/NzoCjOXDMQO/1QP4dR
4so8TBVw1Ig2Pb3Hf9+6TanvNrPmgJtDCMCqzCjthkobjPs5aLwL2MmPGoEQ7TGz
i69MkSWXZgiP4lI+B6MKZRBqharMdOfTzdi4RonuRCA42pWcY/XKqituUjwRW+4R
D8mD9GuuXMqjtjUO9K9/6/oH87OV6482Rsmom+wsPE8bhEk1uG6d+PcwNh0pv6jE
EWGGtf6GL2wHqkMxrztIJGmDm3hZMKuPGVKISrt7cS3yKoUK5ZB00dbmGQVQCJpy
XeztqSsvuzQnRq93XvBbpLtgMQytN0nagmeAFe0EDhwIQZVZJWGF8rert+6uxs6r
QEZCj1jWRXkR0RDYxSbEwF3uSuatVDqJgOeeO2u1qpUq4hnr67vYMlbLO+MsS9lg
vmoOgFK2Qc7hUxYl+L7xtQbFkgGqKmVH5OrQrUm2Kra5Ape5WYTchBUZdgEkszWq
nGKseo6+uLHOwzqcMkt1d3Lt+hTUKSyAYT/jkvq1ujv6+Bf5S/eXE5BA6UyYzrGA
uaWtaoMMe30ldezEbqPRPCQlRchf6xfHavVQ+IwSLvEVz/PXj7+/biMdwhCZYzFQ
7xCu/08d+SXP3SYwCx2p+x1xw4TqtbB2kv7YO2WwkqQWRpBnhjlUKu4pfJTuzGPr
6A8IH5b9YhhOHkNclaR+n7SfYBO8M5HJSDSqogkvaICGCN+rTadNQdxiAvF6Uv2g
RS0MoTDLquNEzlnRxQidT1Bvfxg1hMeDQAZD1ifvZ5iB0yM5/WU5iFgr2VWA8doa
3eBlvavBUOk5T2lL9ROXsOpE0vDYtIQ17DRjfPNiXG+eVL8cNf4alH4+XognXw28
CNeifhEG9R/Wl0SRI5fHvTCSQumFhxtVqcEMW7CQ0pOHGRmXtBPra3f7KkIOKeW7
+2a+ekWmqiBJ+E3VEItAKeA5ntzLzH5c3ItEbdoUnVdW5w0Pd58PqOEwr/hEwRjD
WvfxV9ifw/Yh+QDS/C8pSY8AvIxAzskTVF8CvTlu9reghytZ+fp3QHtkiiLejMlW
O5VAqR11HTdaWQgx/L1O2+dGwrbY/faqeK5cy00UFRtAE7EptCfqZgzIYLcmvGBF
waFAbU3e8jykbNK+Z4UJf327Yg7iUgy11df9rC/H4GGfbtNEg99u4aNhPv4m++7c
5amR/A2H6jY2xJGzqDz3CS8RF7soxMxnXkW1GI9I1HMm3nQuJypkMq1DWdajeYsS
W89OgPQEeq+1h81fIH6dH7/mouWNb1ev5djZ+B+b8g6bufwrEmHjghJbcKDodwMn
ajplU5E2Z0D4AVdx0TqpM4nzGFWT2jy+nWQ6ne05hJLET98dr6suvNQFe7cEwKe8
KLMNPQpLM2F1qDlyZUScKtTwfJyiNVcSsbeGJFe6AyVt5eCtgkxMb7Sw25K+/tIp
fSN9lyjKuJ3erMWkQAVN14b9y3FVTkzocSS1+mMMHzuNyvi3BIk6x96H9WBxdn6u
Rx9XUqCTvGCMpvIVb+ZaruoqHgra50xR5+RkiJCriESThrkQT5saPm7tMKABuEGh
MiO4ZDsb/sVYAkxtI0pGdXFiArcM0UA4WXC1iPJmMjxshZrAu6WnPFbAfiy6ZNMS
tdmHHwKtPQK9tiSa7dk9K4pF0NbUGa9PSX45Gk6hqfWyAxYlSw/ceLRjWcWdjcnM
eD5nQU414VwoJQY1FKRwZToG0YGaEQjaIDVWB7h4c/reKJkky0FolV1t0mNbiJF3
nFvj4SN+AbL70xIVAqzvpHSvaBwKG1wC1af33AB/4K9rapWwE06IaBQwAYoXLf6O
S4KfzEQ1W7b3RE9vDERgf8l1UVJ7yp0EBRCPjzBX3+8ctYA7596wFhxpocQwXKzj
rtdNd/8CD2saYS4xOPzlpMWS6662VdxcrObwUosKMS7pHmWHfPDWceKWbvHnjBU0
Z91RaoG6weFlsLeD9Iy/shAJRDgj8f472v9OQjrcABYdpHc6ifyBwYRpFYRREN5I
NcYPMl6xd87NyDciIS4wn7CmatE/K6XhLadn7QLt9vM7bdL1hwadDOaVMgMrzaNo
2BAgpoGw47wjYXYNZhgxaKxYMqllFgP2CI08I0nnDUMGJCc5BcurpPVUWHyIRSEt
cJz1WfYzO/eYM7DOjwDE/JU72wbZnmqFBGivqTTvQHjh/ToHTPoYiH0u/1R0HKz4
PI+lAvET1CpYZ7tBySB+dqc+eGBuygrT/Tqj9/YB6yJU5F+HoDVPLdE9Nw+4beUH
4XEdK9FJ/pL9KaZDfTtlm/UUoTTY0m7y910XpjUXJ2Tz2RqTDK/PGnc+6neec0XZ
z1wi59Hu4Zzkspm2WfLI689jlbS9E3tDuUvEfToYAMqYaDT4i+CjqH4Ta58QLkkO
xJqfiV4rHdtwFzZSM2ounEJZxui75VTuMbon1oOfCqF2si255KQv77dQFer/Hahl
cwlKyld/qOv0nrc0qT5/XoPo0p9WmI5yiU9QpKM5cICTdqIUQ7N0JryUnfQ/0r65
Dg3aMLKC/LFDzkLmsee7s5SmGHwa7xdgWGW3OnapPrldTI0tv4p+BWukgDseV2vg
a5pE2/fP25DGp1mBQ04IQY/28Qk/qXcyUfx7T/v0ilZxiYOznntVL+Z0JbLZd2pU
KcZlCEp5D1RYauYW4gntMo7F8ooBguKgCsWGnW30IOZ9GN27PDn39GNTU+XUOWPP
/4xjkhq1L+/VFA7y4KlalivapusgAdxe6y05ljTmGM/KVfbWAcQrdOtf4/7wxoOq
3Wey/X+RhRcPKzyrUEyoF/oM65fulDC3rjuMwmfs37U0pLOadzGEGWSbIWKVxvyU
34k7H6cgWielahq5S/W+aixEahnmkArD7HK1j9UoMn37UUFKe3sgy119dAZDVp30
d1NAvj4tM4NOLhBk8JMyIuB5jUNdhV6mQDk9uY6QfGN+cuIzQrGt66XOtJE1MSMl
OuURHbvuY11Cz7h8VgCZ2sG14/XFh+BVbbIKiS5FICCaBtBNgcMZwWbIMyU5F5ps
A0utPWRBWr7nJQM2kFwjstIEqCm6uf1ZIMm75SaF7VYKQeY4EaIK30c7ws92JO5z
QOA4FNJBfrKQmuRIMq1lpQnMk0NVRrwQWvRd/pyG/E+6qU38dOL2xUal0ggS+hQG
Bo1pW8mLDXqaC17e9gbhmnt838bUbhFkQZXM54ghfRrKCrW52QsWHeVAn7t4LfpH
nDmWpG7eU5VYkFI7KaBd4wPhy387nSLO7WT8vTP1CXDHd8rDMEKEvCiJkd+9wCLN
4UTww+FsBgVqKpl6UcgS7q+shLBJ0+K6PaR8ElYO7yS1EesrOAyQmgWb3NiP6BIX
NJv1+WjJssJIms6pGwqgfjZi4yKu0iXJjjz0vGXD8TbFvraVDHplZPDJ4ys+DvaQ
4oTsXhh22r25Lm9zRjabj70xviMDvRmbVJkfVGZW7kR+WN8GtGZrVAzCRR++tQKI
75DUqOPBdVHbDT606jCKIIGu1lEu21VHNmxGrdJ/cfFKS3XGkSGBfytKMDXq+Yq+
BPO0rAmpw6ImC3skvUIopT1BlLSg74/h8WdNOL1CmOuQ98cacJFI2yxQ9dpN6eLE
5VPcilQz0iLC2tbsP9zWPdL5mg2mGj6l+hlcTKlpGm8uM9ZaJhr5y+uh9zWFZkfm
zS3theCKk4M77FrD7FjfBXspFGIBSzdTf/E/2/uq7u14hspZmRj1OLV6no05XbP/
jikJf2OwjcThW71FnHUVIazKbSeZDv1kmOkvAWxSzRmhjKb5QKqozMgBeadlDEOW
AFbLbgJzNSYHY7H83oZtpJdVSu1dSonOQjyUP0xg6c4GIvYOyte2vOk5VTmk5wTY
0efGWb6R7TWRJkKJs0awpJ70WZWpgmY02CfBvhYM4XrB6QH+ULRQJOGxib97pImK
zsNlVFrhpO2cAY2EokPoFCcVYtUPwALQFHZl6GlKGyP+1XGid6L5yvxNFb+OPRPC
NSi32TSeAag8PNT7806GAWKQ7xtuIINgJBrbMkTKLQkq0NFyoFoSIYPX0OuzEQRj
x313Gn9i8aRtoyvIXCNlSNC+RJ6OZ9L0swq7kuhIg0X3VHzabx4u470f8XnjXm8A
wiA14RIVYEBbgdXiY30SRoV8XYL7NbpIID675hOrR9/dnYnQvhcUN60DTZvt3Ai7
ljpzvTP8bxOCT8dPfxEhq1DWT1mbSLtStz51LLEtU6Q7VSZzUkhJt8h+b4TqRTcR
whPm9311ZQ3SX4Z8v7bdEAAbEQAdovUdqjtCdFRVOid3yWR4OeVufHWW9hmLAOm/
d6lAyVPfdmkhx0txYNujWDgFl4VGXhjE7+dtxlI1oWkjCJxu6v/YzaJVyFwqCGlU
4uosptQY9ovF4NgZa7tyXmezWnTSWK9b9P20jJObXByqrcY7j1+DJNmZmIIy8un/
i4UXxcnlQ5OIVJgH9djIQvkQeCkimu9MXLbk8sJBeqJz6rMu/tigzkSir4LZQpGN
R90CC3r710Gm9pYlgJpeIuEdyyhRqR1cLHQBKhAh0sNmLQckrLV/QVoD+wWzkFUE
ylR+cXTioG10e4h2FB0nsV0ROK8YyqduY9yPlMvtZA7q4k9N1cM7IeDLbARMOU8W
lPi8jiCw0VcBeAFvXdZVXCOcMsW5psIAfozkIMzsM8a9e4SPSD7VOeaRwI9RD65Q
Jwb9UDLb32hNaXtz4nPBAeoSYsCdEyDBALbZIxCu3giYewMOGRXA6Fi/RR+wyNKT
2eV/WViRjoPIwZGFsHSm0JPeb1HBKvX4tjCXHffcA1cPEiig9M97YnOJY8cgu3Tt
N4vSb5HMFSNlKtGVkxu5nGVKVX04Va1/sPJUIo2oVptKuHMqickthl+46MgAPUfp
dywmnJkKkSMQMGopYWWBAGKhFNdtf9d/WTFbf90yckRtixmh/E+o4i8qijwWbU5v
1/2Xj6InMl/wBOhFxlhPKqjP0pLVpDgrPdv4dAPHAredL2Jceakj8NdCYhxlVZDd
RVOlMdz9ml4VwSlliOj9FlVDYh2I91XoHwVx3OOWpOoCfFzBKe1qlgRDcI3FoE1/
fXIj72hQbZ6sjUK5uEZE52ZY240Gzt7zshQMf7VrxMtgQjUU1cpGRvVc9LCcCaWP
xu1QjVbbdMWSHDAltTVDd3jNTfI8VKkW4A3Sxh8dKf7S0Z40nFG8UPftW1qRvWOF
aaPxuIIslAOueQZOq1g6TLpr0ZlMZq3XqrFF2YH1NC4ozChEKeCH7Riflto3W8kD
YDJ8Lh6LLjAKy19Q4/CTjWGhpdByaqPlyc/9vvpk81sG8OtKgEi73DX0BbWS084b
i93LDg9JUKXsJpvO/t646cOWZa9CPKOr5eUhkmr7dv3KzDETD9/p9fWJV4diiPvl
lHG8rCiUcMsF9ECe5+OTJcexdoX19fwo50H7ZAIBBWuywMpERpQOEso5WqgrVnHw
5VL+eu7oapgsCetJgox3V46XvEWN/FNOi8QVhbqTJaSxFbx1sFXxvQ+amzl2iEYS
v+CupfW/oEqOb7rVUcKXIVslkps25OG1bAW82uHPh3uF87GgWIytWzbcEqBhAkmO
TcVxwMwrST1yHT9yZGlQIVK9+34OtQOJSaoAm6zOH6FyAMBUwZMlq+6DAfirYhjM
l97MbeC99AvMVEY99NFEu+06t4nOEXis7ZRxgKJemyn6S0ishlPvcZk9rFojo1a8
T8n/c7U2rsczCHqYvYBrrpi7c+HYtTVqsF4SEiiibgnOmV8FKCrXjFotpTMeqbW0
XcU0MCSqjCvnRopPTZQ7xbLMO8hfU4OZ30so12uXvPZL6B4REmzAHCECOw7mCP7s
wDXqJ7UZnalLvgIo0OPHmMTCBxxn+NJt3Jo9KkmuZeuLAGK2pS81VCfIy570oTTI
shTPjtnIYo+9SbJoIefJT5Ni0WVjOb2rbxIBnmVfq98qyU6DE2BaJAsgU5Qb+ygW
ZoX0s7Ae+0Th52UD6Vv6TvB/yp1dFIuAR2YsXpyb+QzaqWEF03w+/CLGpxP2aud8
jtDjdRskvKmxqxe7OTS6qKqiIsVxqGeyOdMInaOosbbuTl5ggJ28rFreWfAYLTtL
dcpw4MO2lf6kiCcyHX6Mo8oQArxGNpVklvxyRmfHNS6/hsiQBQMZud25XXYAs4FN
mgdwS8sDHdnoAlt53+1QikngAMdzYgs5S46cVEj6Inpcgd5//So2RbPi4HevK2R3
+ERwcoKuUrk6MWH2DEEjo8p3CC0YUBSWUdGUnRIoHrXSCnjUF1SqIJFrJhv/9b+B
+4DqNQK6daobYmNAat7qMWjkFTuzAL7BoAyR25ztfiar6AyZh2ZpQwR6FhsRqodd
ZOMDmFshdtaro+ZpGRRwf1t7F9uvUQAq7YOmHJ7xWpc2hVneKzzDErBc2ZRfNb6S
zeiAlxkIravuH8pVtp6UK+ckImFUzdOd+34rHeflWrOfQ0zA3KV8H5e9+bHDAsYZ
rbAg08vt64WH1vROLQa6wdyiB7WoBaUKbfLS9Q0U0fnt5Tf6Fh7InJsL23zDKeh0
jD1pZbxXVSZLJ0W0xV3T5ns4gPXFBZoVqI1sXZmiVaJLVeEGOLa2Nq5LkyA6pbl6
6ChvXDZlGged2FMe4RkTU9JaOWYc0P4a0CPLuZelzqVu+Yb+MioWEK7qvcN4twsy
3wNY+jnojnMMvknBjfSSjroQNTfJzMpkP5fCiXvKRKDmrwktHAWb3peQ/HeWKjTz
KV6A/YzlqphPODRcB4UyCbjKM5N7dBXtyrsiuZQxdQb80Ttw+kewzHs+1uyj3/U/
aKW0X3uG686FnlY97Ml2srn70tYkxnCZ1isiLrqilD7IfoUy6rFHaY4vAeDQk1Kt
EiJUKSdAOCzadr1iqENuKOqyZ6Ex0PAlggLE+bahYdAp3IY6aNFgHzSNGEKE2AnY
DrS4k/MelBpa2bpwEHu9hFDV4c2RDCnPvO2+6C/hY2FCQwCb759pbiis6g8oyJBz
whHPjxcNA+k3lwt/GFA15tSnaG4IVLBYKCz+WuYzhUCLagWwwPJtgJ0xYUHDgS4P
mVAZ7vMhwda6SLA+yom/zU0HINfohjvMlbNhanUQYElnWeHc598C8ZSuG79up4Es
qaIbjlbF3V7PQAzW/JWOdHjjSz/gYFV3i2+ByTOxeAZ0pjDOzQct9biVmEqYu4dL
wXhIK6bxRYnpYY9SoeITdNxR/xiqo8G6BdGWZtIA1ggL3wLyF8tPpqXyAaFAAa6s
WgQHcrRh6Pa2x6tsU33r5QxtFDGXPGGgom+mb7FIGrW5/eL6EIEe/G0gbnNvkNPa
QRs9zpC8EqiCZf+Nrr1NBRNlk6lY/UkmaLYNYxhoznL+kXM3MYrtZVwCiTByeQYO
SmXtobGlGqKgAG6ivjs6DZ0OaGNIapyMM9uePF1P8yd76rwscagPBJZi0I7Kvwik
x0R9IYJGJfJ1XvppEJ5qTtwrLVL5otz3swQm71HexlRUIIPqds7A5b6iWMhXMBk2
qqsksKMWznpvQEk4EFHolr+edLWV4wXEPlARWXKtNAkJ302lscAamTl9gN7krq+h
oRU3iAVbZ0Nt4CBbm45r6d6leRB1SHToq3dd8hL9g/eSHJZ8e/jMyELHngNKQ67o
cRsilArPf8BZvlfcYbVtuAz+yDfqJumjTbXjslvoIcLrRXUv5a72pJyX/TYWI7Mz
0n1Pcp7dT0H3oDlkAuVc45l09c6WL9O0LvM9k70t58s4lhIbh6qZ+EQPLehgVfor
Ttn8Yn5dVueAwHsxaLPa8WKsDniEOD0JBphflrtm0DAN/TZuo/2NT2N4+IwnJZrE
V7CVVWxyZpDWbb7RVK7agRdCh3sIh41+8Eq7BejLKudKAwFRU6Bm+LNobfAwaE+s
5VknLOhHEhG8g+pkMsAcp1p1MPF33rcS4+NlxQSzOXWonm9gJ2UIvalEIVVOVWWB
k+JuTKaTqUIrLr00HUqiXqYMSkc0JWR0K5PPqKLfFIElslr8byA5CLYKOa69Q5WE
Jh1jYGxlXyN5F0ubMwxu4MfEAq7tTa5z9b+dWSt9PaLZPwRGgDJUgkekXwwMCblK
rAbrEQ+0VOpO4nsD68jBMJOEp4cD76umER2XUhvDNFPBGEzs+fxs30bDpktbzQOS
RZes84csfSsSM27DLd3921wD1GmGIBwh3hU1T257/Mql87pnwlpfchYSE4Ocr5Ii
9H5pG1BOOcdx4bv5ofbsfOxrcNE7AldOu0VOn4WzmyfoCnOtf8VI0rVu3mlyVwgv
Cwsd8ZzD/KnV2AXlyQ9KqV8sXvHGf45HW/w66cW5SlkU4tyndreYxg0c9E0dl45c
123jpbj3R/usCrVo0Pa82+chfsf1dgy4Tv+QvTnQINqrORe6nWDC3pWSfcvONDEM
lu1EYCEol2FDAscK4UCuXbRLGKynJtrcjI/FshZblHSpjpvUc0l5yaSMGGzLcaKI
t1h3VJwpSN15BJREJD+wqHjUjwwCNHxWN1syTuHxfyrFchl65Ou8c39Fxs+WcWbe
l/B0GOPKDjsXWpUpiZf5c1dA/IHqae5SIz+Rn44h2nJtBsskwSEz3M2hJy5Bu/jU
DPBEHXbD+nLW2tT6JsU4cmb8CrsPd+5ZuVtZXky2LJyjj94F9dVi5oVf5raLQQga
y26X0JWLZ2Vu65GElQbwVop6J9nXZrgtSCI0WCiBeTJzy1HEJ9W49uTgsbS+8SHF
997v0jx0/Fptncbf9MgbacgGeKEvzQqnat3rA8c3Rp15aHBjsm4fNr81hEsC3zsY
z8i1zFcOrDTxxuyCIRaag8tB6ZzZ/ykHugbguO3s5QA3xf0608lS0REfuePIFH8m
wf/yk+ubIqU3bW9eoReguMlY9zjb0ZugAc40R/9CrYcUUCVudJy2t2JS0zXMv8D6
at3ae3VTvz0/Se1W3PJSaayNvj3TdZ24St5hrgkH3WyKuLrhrGhzxif3MZFXYLsM
4x1QLXAAyjivfI/dUwI/3/HqW6f9nTlSOm9h8NlwbpscicxJmLd01YCk67WcEB04
qMW4f5IOKspv63p1ZTGwoNBMU/9VRC0VwW6SvfK1ODg2kQLZKh+sqqnf/IK0Ny3q
RvTToHrsAl16idnWIRPjldawW/BAFKUs0zPhCf3xXCO5s/8IuYUK4YTUFeSbtAXD
lg+H1RGNoZxoqSEDCzEYRD6QDNZre8nX4cqxay/YYvT9UJxAScwx5o4/lEyMHPkZ
8DMpqDeKAavVExh3Of5H48ocTL3cFIY5rE8YxK3piQHwBNFbGrZU5ItZyLjGqWUM
A5Fz461q3UEsbkOoKsI9QkhU5N6aUa3UtVFPDnDyuhSaiSFSBd7viDsg0l/Tq9dB
08VZ1UoNEq1+sHFogZSM05g2UEVK/LPBtfmQrAl0sC+9u0EySkl15ThCyRVLQIfQ
h71wTFxWNqcPwEuFI6VV3QggZ+C0NBtnlQMsMv3qyDDwne9lOm4cln3xjovL6vgo
HCFkF6337rSURsySpg9tLtYRjja1rA9PFvnFG8l+3w+DHYcG4EoTxokXHsD33EW/
74E/H3fGwZUyNk2HYYdMx2eTkGo7dLUA5C+4XU5vWpzSeA1N7kjx+11L47KN+VwJ
0MSgdKO2tddmVzZ/UCe73adKKi5UEcztoSc7mpwD+9nm9Dv+9dxHslQU53LEzAbr
mbVbK+EzNuaD2pvLHzt5ljv/h1WEo3eNHFc+GNsagqeHRwUWVP/jDH5wLhKRS49a
kUyLyqfsO7p4mWOvtGTPTJZLBz3DKXhz0B/Ya9q8nlmf2J4mKFxbnXS032/8ZVMB
fG1+YwPbjFdUWgi/PbFDvpEjidR0MvHxkfBnQg8ODbiBz8RM+v+TGrxMzDdNPlBb
LLiD2rjZUX/UyE5BBCxfAlEJQtBih4+gSascclzvPGG1fN9oiaBNWtsu/bE63x2n
i6ge9i3Eze64IIFr85If6Fkkg6hgM6xn+l51dQaXKJgZtXFEphEpI2cH6nLxPoL5
N9fYxfZPRtK9NGYBrwD0WtyQb1FqAJ9cslDJjLCcAs0E5JyQHNah+sFcqsWUGgHw
cqNDZyBzjN/K4EynaGiuzPbN6MbfYfYPQMDEEVtkEyYUwG1WGuL6jkG9ooVNHY8b
ZZSh2edcbl2ChcAWtlCvBsViFEAufxPuzNHPkObg4ioXB6pyYtq6alkry5R2Ds0f
5w18poe3ObTq9EdK3o/qqgJOl6knaFV/VjzyEgGufONm8S7hMaTOwqY9idZ3kzPk
C1ANoNUp6xgXFicYgLQTNPaYDGyv2KCUUDRPI9NQug1T1CrQKPgNP4mV+mVUgEiH
hfP67l16Hni70s/a7dzZNxokZCOHesLJoShZjMngj7ccjIs+jSlJ+NnpLb5zs21v
lH4WgFgTctswrc2xE0azeV076QmwRk0kY04dMgncqRJct2825U3XkxbN0wrZnFWf
ocDK0V+GD0EFKPiiiRBuCvH1UiDInySd1ExXMqwaPqjpCQOMixcRHAMfKnaOHLty
Bg6KJazdW+2jGQy1YPzss38zWc1qbPWSffUYCeXeCPGcaDa4BpKR0nF5WgA6UEnr
g3ajwHKU8q0Ot4qlhQZJHHOwBXndpEndCNNHx6WdkP3GmTQ0m+SJO37+zA/z4HQZ
Ulylalrk2reCjeO+9zsJrBG5fMqqidBH+X7erRDnu8CVSRp7X6yjMXyu0VY7WhSW
3piFI1p0jVMrx0Kf2mQp627PpxCX+OeYY3ZFFUucv4HAk9vejSoj3qzvMwqXnCCY
n1C5fxgaJB0WV8yHQDSRMwfy7eLzJb6TuJsM8sAfnjdLeeMxZN5CvzpJB4EK4Aor
9XsF4NO8mQAKZy/NV3fhCwEHZD3iOVJqSTYWQPrtaEQ1s0mhNx/sv2WmiU3OHELy
EOEzKZZAtLuJqpPoOGpjiVsasxXE+xL53jlEsx9Y8WqE0DNdoCgUQH0rrerhQtuW
amw9PyDMnWcpwCBgzjt+vBXW1bvda2UoKR/QZn4WrqFuOBYMP77/6LMIgL60m9nr
73LpNYTqSUHLrjHv4vmzy7YGo8ZgTv/z1A/k1bW88uhOlL08Wy39r4gzu7t+qD7/
5QaUYnBTglpg1IxTpHigalL+ekNf8VmIomqUemvaTxkFBVkA2L4TOyC5A7T3Qq/u
cApBpeVyskrE0gzPCP0Pco8nUQDlC8XkLcta4JKccnT6afdkpFv2qf2nWXzlaOLK
3dJ81J2Ubu+KYkkwb5AlE5fFLUGG3h9Dq/QGfyRRtdTRP5MQuE6rkWDYDSrw5IWG
DWMtp0ltR3Ct6n4n/hRg86xN9hZkLwtnWeSMhz88qtiYPAL+xRgy62HLn117KcfO
RBUFy/CLMh27PlnyiwieGlqPbzyFfmbDYS30SE8HC1EFgI8mZB5i2BzScyydRDzv
iWQsAjUsQoPa/ZWmM5KFr+IRT3wmB0viq4ZxG8Zjt+lXL/n1TGo4j/dAfRWvSaTJ
ysXnZVKdUeYT6m7kqcwUM+33LWeeyV3v3H+QoXEYEliBfmV2dT+OtWAC8befqM6K
Nh+xITAbS1QgR283Wm/d6X0YFBQ9Jh3NGMBPKoPShVr3YLcLr136CBDsuy96xUhZ
6YUn3A0jVgCVqUOEDdVmfSnzlf7Dm4QmR8zFgwQ0oOJfulrclDGqAkL1GBgC5/xA
txJ4f/Kx5dWlpqx/6L+yrgs6WJMnO+EnFIY4ImcogrSY30D30yjiZJB0CYbua75D
2dZxwiSZmSvE5hMRZChqTK16YWXlwHSReqvPzuOazqkrRhhBdOQCmTJ+RwE7VIvJ
7w1JMtCohmua922/nLNrWdi6mP3tv3/JgpXbdWp2sUeYyIPcO3Pyrqc1qnKwtqUT
Wp/n5nYuKjyxyiJQJp9oSM8cTRuNXAf2F5pfiNrBiGnLmbkUjP4QtdYCDRZLmCEW
xOVwXhwZQdhUsT2sEAgk+z/fk+Y7A/FLeV5rgv25RHSZInsm0iGAPLXXGvL4rjkf
oZMCxhYI83S1fuCXecOTZjaEyomxt/R/V7FvZTYBgcBQbLi/16dh7fQ8jPHdBJdW
wohELMK4/7a454roMuRdxj7NHBniWeiVX6mE2xSqZ6bWuiq77Tp0tgFQbwnX0Eqe
cSoLAAGNMMdSbFgiBWxueAxdz9qIO96Go1rRB9Vg7c2pnzXcTtQer/ySLSafoPRl
aVfFp5wjNY8fvycjhNqVk5uVFSk2Kis04B9AZL4dwuujsZGvwlrQAKIu8qxkwgNI
NOWzB8QgO2Af2I0QpS4jwUUIA6gYDLMRv37mljOJ5k25rxWnvJibTje3PNnvtPfS
9JOzAUgCJCy55/H3vxMeHZsfV/qDCMMhQylXotkCs2MrrR5doSz5VU65fuMd2rJB
C87ZL6mAKL9mWwL9tBJHEH6ri3X5codwg7krH610GcrGtvLtOBK7jEeLqvBMN4QF
BrtSGjhwIpxu82NlLOTbqiDRuullZPgxcanKP76yFWhWmUoe5ASifDgtVvzIPEA9
dJvj22ByiDFFG3NYKe1PwlvKHQac53mlhpEH5jcz90QoVpPoydwveypGLUGB9PUY
ZeHIIhyojKR8yTrhP25cklhq48rtENf96iIfWuU9lED9FL7GgWa6v4DmD8EkGdiJ
Fdh0JC3H4K207jerwzReFmcvpodE6KW1E1ujdYXrM4V/EYMtqhY19xXrUU9NgBKT
hjIUOCH58xTD0xfUtHZwSvMMe1+0858KwhtoF6dvwhWNulrIzpwGwg8q7ixoPNyV
0fx3KJmxYligo6gr6vHa1lyoOdTSXt5fnPYNO0uyOaGvA45gVSlliSfgMdOCIVDJ
3ZJf+HauS10whaQHrA7cUMb8xLSEYrjtj3OGc91H4z8/qd5wOgCRhp/bcsZaBy3V
ThsHfjEYU1/l/I5v+627L5xSPkIuRBeCDsqu0uTxMJH6BRyO3vcZ4mMPmcmUGCcd
yPCbhisMPVDcgxhb6uph5HNj6UXUeBhrOue8IR889rQUdEn7xyWE8H5qIPPvGkYc
MOZ157ZgumZQZ7RItL0vZDYqkvt9IDgjKq94YlIdu5wRCty0q6faYPEUl9Ykuatb
OVNtiOhS6XJiwr4WAloTia0EGyyJGzoHLCXVrlW4uLCwhwFpESz57EQ/2OVTtBbk
C4jVxzSxI0huVIpKov2I+Tn0SXJPEUNZdXehvBzGsisUvykX2fWMd3/HhSZDX8V0
UujvSPEAUZyHXcmfDu8cUyKedQDgkuqGfWOxRCSU6wT6biCEVK4JZv6+xT1zD+Bx
bhT/C4dbQZo4D4AhBXHRcDqThX+Bschdp+nQOSLUrQZ7VKa/ylYxMPgyp+cn/rfw
l+8+VUJ9AmYq4opzbZ4mBnzJ/dKGQ4xQk5vaNWQhMdS8g/i5wvWj3WDlnGCWs179
guQlSPX5vL5AqfPqdIKBTqVAa2MuhIpht3KKZU84QVVHIXEBb2miwJqhq8S4HJKS
sxmqA2kxRil7jbWwM33u0Vniyq6GEb1A6r9uEHrRm1TFSlt+5Q6yFYWuNfzENFZV
MupDrC9ML4g6uQVyazPz636TbmSV11KKkoFHR6e9URy6tNf9RC6SZXBVOBBLJ1CX
N2CbIK2VN8WbHvINbJUAnx1Itp9rChRs0nl1Ydir13/J2MlCB0NoU8/JRC9JFHcN
PW1wEiGXOwnUO1Dg+WqrDLaoNCWY6A3vYwAQxDqEjyJRscReqCIDGPtvA2xeubeW
4i/gwXxa3uHjP/Ftq8r8XLpoH/tTrJDc00pMc+psgsllkS25ySQhgTNqJ3d7hCrg
cM0i9JXecV8LyEIWvyjpR3OxH9+7M7ypDMpOwRd8rDsTK+0/bD1ARDerZkzraRx/
4UjbVOWaGlXT77H43cpYhQRw4t8nJF4q0SA5NzNs2pbtdjvaRcCTYkZgWVA2HZfz
3jWwlwy9LV+Zrjm/vOAzv8XBN4TG8rfctsiFilPD4mG6FaXdIfbmKKoasKcW7FsI
htT2Cg4CYNJLISAV7WpZ2aVYjQmiabwhe1rRMWxHbeFdjXiHuo1dFFnN9rfAbQG1
dL11IybB/lByYTS+0IzUJbhIHoAsTtyFTDa2yTpsEBNkCF7Mt/fCZ+RMyojOxgzF
RwaVlxfo+RgiCjmtn/f0/GUgHQcAyMC/kmPVzgeJfAx+breCMcYtRublSmZIAzIE
z7Qx7Gi+/YGqilXaSR/Su/9DNw/DOkBXO7MlDMb0IG045ZeHePHuWzdpu+ruD3IS
Ar/y9pNLWurDzKnr3XKAy85L3dT0go/2joAYcdCB+Y6FBLOUbazEzjSw56gDzR06
e4n6wUTtNK7XL8EWsTFbUV3Ak4gmRtVGHGHpo/Rg1IwvlzKTYc92mF/jmuokFXtK
TsDnS7htPEvNl9DFNV6kbpS9SwJS00OJRjhP+K10K33c/ZEgT8phNRjWU/YZs2oy
aHptawlO93AVD37DKAzFfwiu3qCNbg07FdrYPEPcnkhj3c0/dez38GBNAQqKEq2s
KxRjHzSA3D/L9OK37cLmptBOgNRIMnh0m+9esCjBMvOw8RTv7wxhZDIsIoYWKqfw
8HgwfaO7kVNl1K9nRnZfBMsjuLKC05g1SNbbzEBqH/A1dBaHejIxHlNe74gB1nLQ
oVle9H5mmwm5XcDIulMH3iQvHY4IKTEEFKsGIwUGJXiyz6Y5J2Mxq2f5ryX+Ga9B
VkbacogQ9KSQvPb8lTgWD1W00ZI3JUVF0mUlX7v+H7fDDbzGhPXPG3dqDPl7m8Y9
5sE4Y9E3lvUXHifZPJcIIIHdfaDEGweHb3J3b/T3lOtZFY5HLFoLW2PS3HFNMDdH
8RHQAuuC6jP7Wr4DlYkvwPvFHgGo75jFos6qMWMGY3qEGAaAwTFfgAZeKZWJL9b7
PdYfvwCxueQ0fR3oBSeU4PWQm5u3hHqm6MJX0GCVNjHJpc+FoFmFbF9ydwk0GbfY
7QA2Ed7lIU1NeS2P/9mAkDFo1W+BA9sAZDEbqoCES6l1EsyEvGXlJCnoiM0tLU4X
6RBedivGGhAE8lUU0IIqUvcUwOIT7w9FNpntfotwcfqSMUquidHJYCmWGO0wEfbr
jISVGborJB+i5LkKC3ObVogAuPijDrMMhVg1mjghXu2RBcTqoBIdqGxGmB4d343m
jSj5ElFWDPpt38yffH0tNoc2eL0vkgNhwk+Yq/qeiSeXVdqm8RknyNFqfiWjq9zc
6q6MNVvhHOm5FWDxMJtwmthx5pqu5VSZ54fTUvYVmI08XkDu2FZ1cRoii2WJJqD8
6s+WEvuOcvOXlEs6fKeK9f3WZgj5Y0E3STgNLPoxXzixpraKmdTnCVYIRsWoxBSS
7LVGY6YaqSaFhEXywHTV7Dx6yYQiMiOWg9AypkPI2/xjlGPyH6Xe71JEjhQGvIOC
JYiQ58CvNphv6cHZXs96pEQTx5710g8Q53OOuo+P1yrotljMpmm8XM0IpsLgQSki
Q+WxpV4BTIJI5/QcyCJ5/VQXSnPKmLkg++W6Z7EjcSyJYG6dSKUraPETFG6v86+L
f4HEQr5a7PJ0tUr8NWzig77srebNO2sMO33scMg8Bssazo/GWQOtOPH8p38HRURb
eNhhx/4TQN2aJtjyHZpe2ejo6FXYxmf/s44TENpROiwHfiHZc4ovUKFXl1N03GaF
8AmzKeomFx0kqKUrYdPjmM+u798fmX4nL90RJ5jZz7RcWwymuEHESdvq2Mwr3jhU
a/lI+xnp2wa0Aj2V/ybp+Ia2e+ZjSsugIen3TircgMlnrqblV7nAZb4jaBxN2snj
4tnOUBXOYAfuoBlnbHVj4eHxu1QNJmbF6biVYxDst+v/rZ7ivsn5N2wQ6Hssd3q4
KTf+2GVIUdc/bnLeIzHtDpFTfpeRdT11ZJEItX3POteHNJvNrKTSFAtfyYaH1RCu
Q6++ue43PPgqdZ2AeieIlxq5drQy8jsXqXFnkXwzJtVyZZWgBg0BIHwbqwzgJkIy
jZJfShuewNjdBS2bc91DGL9eueen2oMQvkD3nmnMc7d3tr2o3XmhG8Jaeacsvswb
B4grhl55UVSDlDitw+I71xi4eiaQyG0B/PMeFotTeYAkNzocHbcmBrmbRAHQXDzV
Bf8UQsh33vYbWIoQBZK0NC642gXjqXSS8Y07wwm5bT82JUPfcfJhvgMVgTsmy3ro
wgLiMl503StM7QE3ptNXEzz9KvKf4QUREsuTBUIIa54qYHqnlxB6m/jw0s1K6yiz
XrLsfvtldke37AjZV2RdfHJtAxXeEwe3IarrILBoa298kj7AJAz2LvLMxXJMmhMZ
BslHJryIsSmfFDNB4obqrtKzszlNpguvwNHzl8n7IqujwfINxXoBZXSoNgrtkhW+
WaT3ZtWoJBayOEOwPCEhqB6X7Pm+ovnUxEjRE3weyCHymLU3A1prwIKjv/iRwiWS
pPRSG/2OcPcPQb4CVC5h2s61/Qk1SvgpI6WanLvNbUXQWzWr2NjznUqaXZpedKyS
rRGQ5zuUduXxWVOAW9khGZsIz7iG9HAjZJ8VNaipUtaFArRS4+fnwkIHTlaAoWNb
tG/Nry3KA/DIKF66F/Aim6n1OgqILD3yTAg4sc60EhJWaVwek94kNVlSdgi05WF1
HpS2SZ6NM4ivq09LUCEyNckeT6ml9Oi3NkyH0RPhlh4P9dmc8+bCuSDPmZ+8YmV0
nMSAgrzfBmXooSzHXwWXBzC9iRBfCjRZ5VXow/reNHBi4G7TCf0IoQVynoOT8utM
X94XPomZkcrvgv0CNHYsFoZDUbVb2qTSSGXoWZyWB7nBGu9QSbk+N91S0IhllJiD
1UaL+uErqhChU7DHivilyq27fq261bLacUpwXcxLma9DyffdxP75WbxQvzC9Fz97
EqNRDVkG6s3mYaocL2hZQMoRCP8ptJKCC8XTdnahTrAPhP2kimg7j0klzKK0FSox
bqGiF9AODrevx5Jrug8vvI1Uom8NivgJVD7ozJXR4sv07rReAS5ba7QD1Mnbk5aj
WT/UlOhFYQvbiA/8prLchAXIs+8fjjR43iOgjja72rOoDpBOI+Z3xTkYHGpxqCOU
5WXfYc2lnQOUMVtn1zdqvR2tbN/x4ezhz2L+sBQjyXFjKfLDuM4dh/vPg4Fo44EL
IefX6p6rlsSQwxmlKkRdjqmx9TQ23RCyNCx7ay107Qn+g1AkHfWxe9BJXnnqdqtE
3eySlwvZN4mWqJcYEg4GYTVAuaLu9dV0lbDq+XwuTVQOKuIg9G1wO0KP+s81f/nf
7XxRS+o8gwmOiTjGzSepdtxP3gvDtCt752VDbQHFg2lY3sTTbMJ/S2276aZq2nWE
zDm+3Xx0B9imHxOIw7h61iZulisdXLJxQQ+/W2GXNzadVjy7EIsLotkgNrS7I1wB
dQi62ofK/yW7uaUKXX5fHHqMQs4HfMIABX676/b1b4dj4UOYqlcvTJrmjQycUc8G
2LbDnfFYpUWbOyFqCLoFCQ5ld4eNOLPMVrN1MrA0iQrwwScIiyLbU13zAe5emTPK
VpcPdE73IgGfRVg9EnE04JS6bOOrlJw9pJlWW86/fAYRt1wW2bv0a8GwEz+0S7m0
Clhdrt2oeRqu6rdncEzwqDBLlxgc5lt1Fa+ltoGaAOo+XRYwjl8uyx8FeTqgf8mJ
nXl0pQdWo8N2zFxRGt3T3FVgXygOpIjpqREa5XahR8pf0twdc0xKAvXYPLa3pAMq
dBExVwbzzs7OJn9y/y8T+U0iylGqn3CaeVYaYppiPbtJTXvYE+IyH8VbWyxN6el2
wMLdjMFhWmlyqbZuiJm0hHywURojqGCkLDTEbDzEGxTEPu0B8IwcvpPevkZUowL/
l3scbkIQD6RjEO0n2HgijwIer4aUhhazjumRkqyn7TSiv9Kbg4mMqpTTDg8uTN/e
QANVHjzt24b7ggqLLUNlaPtb5z66WnWG6/jW5/NmW7tYQEl0qY8H7XT3+Yv9p1y1
tMrRdsnmLHI8BCPcXhgNOexZWXr92XZWrwTYuT7mz384HiTuyxVjfaCEvP+Cw6hh
RlHY5nUmFYmdCHlbE8Zuvce5dkGv6uiSWsFhKFXsGZEHPGX5vVa3B39O6me1aJ45
6HlYIp7uL0/Dj+4BOxnfkerZbUoMmHxpexpKxtEHbuXPCGBbLNoeV8h+Q/ZFzLA8
PUFhjNN9swsAparFhWQDd1nRLgHLtfRyGIxV1pGaLo3owdTZsosWZA2bJSQjH/s/
OMlSaWaG5Puv0ayyEYGvrDj4zGos7qkwf0bEw2jn5Hz4MjovpgGIsgKr/ZK7/lU1
9cOoPETFr9QoO6f2oM9wLmAmtNmxK3HD1nAVLPI1U08CnoqLnW7yvyrZLK6Rtvao
rxheiZ4cu2JH8XJsPTrGlvno/XIS+5RMk5DDUwfzLVi9tkArSnX0u6JeRpIStw02
Yii6jUTcINYLwfG6kLcUE3jmNm5czw25Ms665vlkr/d7QQmLaBbQr98cAE9k3xQE
l6LT2meG4rmKgHND5H7oq4YXuNUTlVzs50AQhjO+FD6MlswkjQTiilkWHVjQlloK
y8R1bZY7/WdF2V/VU6GQaD0SjpQuZjUPKasYPJXBlNf073VHVuoPebQZnEe1CMwc
mufAknzMcQkpa9HQHOYfo6GaMoXdy9j/Flc7Hj8WNndug3G5wjxNVgmSha7MzmDa
RsB7ghOO8fg2L+d7ZjHpv2DP4kILtBE0MnB71oI1SwuKZjSMkW6yKFm2dGNhXNRx
u1RFMONXs9IQwVfg0nn/T4JsCK7xtgWGMvdnGq9U1+BeN1VMbDXgYDFh2Z8m1ySk
GklcnA8xmLtxFWENI9Bep9AiXNAN/E7w8UHsgpHil2cQ0p90G2hCqzzrdIoUFRMe
zDD4bFjPKOmwJoA9XIMprQBti5cQG3tMeSGAgGvBEaQDS8sIL1iJcYvuGTmrt82o
i0yr1aneyXlyG3HmA6eY0eLrmpxFoFiE2MgA8ryhvkLoFYYEmOUaaIn51FWAGbSp
UKPqEWpiQhZNoUCktXYlkFiBxnlBRiuoggz1WNLVhrf5CvJGnv3sF40nga1JrYMT
9RXqLNHF8BRlyC5pzojV3SL26daavIrFUzFbp3zE2AoqWqIL761YD3OkfT9Q8oM/
jmdf0AkhlB9fcDdSso3GbhQ9FlTVeOxc/ZNxmj6k4Xc/9tMT9AY0YTVyEvISLD5j
2EohPaYIddI1sOq11b1AZhgxY27CBsxWLFb4yQUmYeNZu6YETJkPKDKnhxPV5oE6
fYuC8EcbbssOnm+J4DWjKEAsPCi6S6Wqr+dGHOwN21oJOjonGt7p0xStVN7Kk3kZ
oNgWhnyzObT3Tf1BJCz9wLH/UZiDdnFTiOoAcq3mz0MfZ9O9fjbKN1kYj8ZVkcke
48ac8BKM+GTgEEyLgNFprbqryjKu7WHB2HmuFOWt39FmihjmNoy8xVZRxHsQWRe+
tAqLIT/FQdC50+c1/yCjcBPGHsuzpIwc9bgUzjQGKiSsZDfO1KKOxvzaS3WQPxAj
BTe/RS3AQmx2k9GKNGu+sOzx1KCacYU1q93/dR0S6u+YWd+HSIe3TFUe4WY7xJZ6
qCySX+0n33LKmc8WH1taA5SMBn2KUWWKhPUaEgYdBawrGYNSupeZCujrOkXxfOcD
yOZFV57Wq3V5QA2EkoWKgFCjFBmWBghxF7fGpVzJEB43FuSBVD47aQb2jY7jMCvZ
+H/iRXNFjIxAhVKbA6EhvAB128yR2/PBYKBCirLGuPNnZW91z2SijHoa61lWLGBQ
xEEA/iB0yKUOb32iF/o41WKTVH6gqvKliz32nszKjK9ZWWzVgEF8vTKm5tmWXUrb
KTLOJUsiH0dut/aSvkHYSXmMr4HBFtDCwRyZl2Fh+VFzRityR3z5JU5TlJL53k5J
WlayZfLODMh+Cmf3zkVJjX7PQO7QPogpjykA2TmU0jT8LEa3IxgRz8MBND68RIuS
XZeFrGKwMVNrcmZIGDPNSrzPBeRbAHzWvbZZV3FS0PIpxaqNfeVtCGV+nDmanPTR
o+gxIhUwQhcG4rRsk1euzse9BO1BdKE8kjSbafWFrLJEjVhvAEuTWHLoZUCb0Ss3
aZy7ptUA25JJxiiZwGcRBy6imhPux/wLCskc8mJ8bbUeg2A119gmKRTtgMaI5MU7
159OrpVmDjf0Pv3r9T5UNqvJUdSrzyw2T0f6yr+xJWIbjEzmXDtDY3d0gzUen0aZ
PUnpiNSbJKtjIy6n6r8MclHw8ESI1UxEN+o90K1tIAhgN+cdQn+ebFe91oMIeqPA
qtFINukLL7yVkrNUdMDf+tULD0KcwAr8SaEqaSDophsITSyCq1lC/CuOQryUEM6E
0mQG5gs8PEb3XJHP/sh4SnVelQ7T74t/RA1EBDKnkL4BL00FU5+SKCsfh5ZkyZvS
wYMyPFMOlfJaIdEPkbZzXdhP4HCyGu48PPUgD9VTQFjD4w6nc2cxYBsBMnN5mR8l
RB3ABJ2YLxSL07/SmUa5W48jYY+/tRauUZi72ak+mLD6z06q83IkvT9RxW7NbLgX
ztvg8fcLyQj5QjOiFAVwDb/gErgcAm2xTAz1/GUdsMp5tKjDZQ8ew7yrei3hUpIl
fhzA00bnsXGiP4i8DM4l3kXLT/LguypV0PEt3fdtAgJKENts6N2Qksqa86UqA/o0
WWFW1m/4JoiQMbf4CxrvWIgA4kgfTlI7fM7njRETFphHn1K246NyE0pUJ+2GNpWJ
QtbqYSHbggO2V+DXJ0sqjYb7tNFMylGJjj78FZAzrQwbpZ9oPvTO4/w/pt6YnQSb
D+gkhCSE35qaOntOkrsBA6D0DT0zSESQ7TjG+vqQH3rexIyZq9U9HH4flAwqaFD4
/Cb6e3LiThrNOb87wIA6zDFfZ+5G+f+qWw10j+qikj5JTYSTMKTG0vL2Kiyh5tab
EAqSc1bni2xnn54EEHCWAo+x1xiM9jRI0P1TmffqJbnC/jTF5HQupTbrqkhDpHeS
rjbgcWhJpKKSFX4DPuiZhtUDQAAjWRqm3ISMX3gRwGn2UPQvyLdfX1zJlGtI3K5r
I6F4mhPh9fSEhxXFsg/bBW99SQ28XLKhyNxGbA3HzrZ0JgLBwV/XHamqFqfgHtNg
NUVkVPHAhuCfwMdo2peDDKP/G0S3ngPUiMMOdP8u6RDGhYIcmKPbzRyZbvR6tASW
KA26ZfuO5w+Yb5JP4oWw5niExavHNLLk+lHsE8Cl7Hu7oX3wH1Hr39ZEIExAGwFX
ENXQtcrYY2u3arJyUD86PGFpw/52tOc1uoJEn1fgE+bzvW1lh5Oy0cuZjfi34z76
gps1sbGdF8SQ8VnEUL0lGcOAkwrP9yaA4QhcTmFSC3XMsS7ECK4LVFWVVQaX0Fqb
d5xEOQ/erZ5KjNxeMN9csh2n56lFh8WrVAJ2Ga6Ny2V2wMwKnuBaqZipr4Um5CNo
i7y7q3JB1FiypVRMReSv+ENGRmjIO5kQ2zvkPjtu0b7DokMWSPca2UQqFw6ZDZPZ
jhuL1hoUNDHFrYR0hWsozJVsyL78jzhiwsCNpNwQgCxKLltUxwKlznH3FtCCJoVn
CzJHUVS8q0kEwl4QfAUIip+yZx5Gw3mm0AJALMBbYD3/MFs0mxA3O6U+Qj79KuPG
yJLyNnyIZ0XUIJ7rY3m+hcIWCTpaPH9mMXlgTPuZW0udtO93FndkQZXF/GQfET9K
GXJqskSh3pK4CgEdc4XWp2Se3qMFA8vTeKawhito+RMRNWWe5Az8JNxG6W9AZyd6
Hscpf/ijCIbgr4zvmzRGFaithi5wRjMTZpzEKYJ0a/hK+ocfETjzfoCBV07iEXIJ
4/M4y/uq8KgHGV14yLR7RyTlXFMxK3jIti8/MHCLyHUjmI5p/9JTzmixy5rAj6Or
6LhAdx2pSzFcIAfIYTb6IaAS8dF4P1igUN/sxfN0ZzvufUYppUBiW/gCGpXfazqe
FH/lu0N8u0m5KymivL9R3I0QuKxZmB7gxSYvPK55hAoH1incxyexGTks3FiZ2t+v
5L2IPbMKBCBEBiZPcm4nZJnS+SB5K6OmntixJwDUASopCyjStzYq6BMCzmku+fEH
3fdo2rSFg6BtbcVQhrJC/XQNY7lCxLGSarhhZlHCHrd4SUbsOkPR56FC5aIFxvG8
LdHOHX1bYPwrLANxUzV/wsd6TVTy+OXvSGG4HO6KLKMmlDDjABAFChwafJNQTA+U
DTgbo8B0EwGydA3ahc2TWdL+ZqAip1C2xl1DdQww+5OHIQzbWNxoKa1NSA1MYJTg
0HOdCZtIGbvfb/G2T5iPnTTXkBIbkEEG9bvAJMJpk24J5YLU4v1ztLkETHJYuUKW
OofUbH4QEBRjMrB6ngd9CNQstEJICDD2B+VQ4bqQDXhA/I6npmvZMsbyxmQOxdhd
3r2ytwWFkkgKAQwDaUAE4TIFFfJo1rdyW/sNvpR3oD9iGM44WKDAucpBOTevipqh
VxtghiCD9BKmfN2gkpj7k5Hip6t6HBNQIZQViN21i68I4KprSfaSocwNMd+KEf2q
mcqR4B6FqpsVeO9xjI/NjF0M5i2Ytzpi9RPyCFsoFJV27lbtkAK2hMp5slSWYA+r
UDc9TlK0STq7/73jRKnoUy0YSKiDYcPggvnC8bMwv5nLGSR1nnULOog1oxCoNfQN
nSg4ZVhaBb2o6SPfvlxNh6+Pbv+GPIwRgO191EXSKz/T50sA33M86tFHYwaTogFd
SFrMhUdnHReELMz+2SKBZ3cWXi1EA/5RLCp19qbIRNAVDv5waPfO61JxZ+JB+kKV
fnErxCwSQu4HcookAOwsz8rivHdJAloPFC+HsRkNpimhRpcX5RYd6Dw62q/HUGSF
kRCvXA/0KPae9EWem+TOStjOLH86jS77GEJi/kL/9WNIVyrsYKsk72Rcdb8HA0vx
cQ38hI/9XwAHw7kMbx+uFSw9seuFUFkxEYKPzH4HGffvYSqpPPXkXn95AfiunRFd
MILtnxU5zOVDSGNqQxNm6FvdINtxBKlsPsO7yWzYc0axNFRKDU4Q8IKyuUhovKpD
/4NttiwAnXCKYlruc3bmnRgGl5n9mwbCmyewBmmzepGoo7QHcAPCWt1xhtVwOR/K
7oGXls0mS8R46ni5DTNH7aaqX75P7qDRRXVC+uzEbvxkIxdWQib51exly88Iub/L
XjFaKMhbz0bG3gyCPI5HGuhgIrMxP3xGXkQvVNbuSQ2xfdIyCtFr8NwNDdl+L2HN
yRld02oovmZeVyaw7rRgkbupAJ3LqgDFX8nHc/EeQij/mKNgv4L+4rBY3DTSaMns
IMu2mWAD0oQRiD/f9c8tPC2ADBeTvhYNAcPwioCoA5WCNtdZMYlkaoHnkQY69UK/
MRdxGiBNHWxwP45zymp9k+54/6xJaE3fgR27xCJK1Sia0UmMwpyWVACM8VTOBpF8
ZAAR9yvqOBvzGM47wAlOBfhq4QxiSof4Zoo8gOcHttQCoNm60xR2yxn5D19vUIYo
zBQVANQkeZDQdy/ohZk+1kBmapxtXP0g4ujTcDVplMboMQFzHSkXC93D0vhU3a8K
d5panM431D3xqjGicBO8EK98mf+z0BLMVLzOmo5G3dCy+r715zdB5sGv8ki+2U9X
vecxCHBOECn3jvd+Jbpl1B79SMdPy9ANvnJr6wGXPzzF8Vl7wodZfrhRKm2AxwZL
CibPjkjZq+Qa/+qwfUEXkwKTvt7wIEp8Ckgtbhe315/JoZxlf/wMzbUm18MhQjdW
jtZ66/iOaqATqKme1JKop1ThJ6B8ZbJ/muEVaO+Xh05/uKTcxm+sKrZ1Bl4p8hXS
mR0OGC8+QGxKl1eZ/toeaXN3fe515ccrYzgDOfOG8bBnretyOw5LlWBffH4rmeSD
8dHQS1+lmP2nfdZR+Wb7ilDTN4xx2sGCshUt0MJbs/5ullqcrw+BAM4vjTUOQO5F
9vMzfr2M0lOEO5XGVtjQ9Vt2jpPLcM+gP8n+Iyv7wdfz0daITvVlC03fiBDyPB7B
WJrDq6x3lZzNPrnIzRr1JgX8TM7aXelwTw7B4yeMk1yXxaLqgn+DIQauNkpnJuaz
5l8dbbY9/2xdCarRNIh4aTsWCqph6T6OjbtdNY9BYNMfLL+giUoTRy/u++LE1H2/
i7iGyASkl9YmVAK0K82e5Z/M3spD6ACagQb3VUD84cns+0h9Acs3RKFllVnDa5eZ
8eK7sM4/bDSo3S7LDXqywbVO5SAM3snL4MiLTl3RAh/SPIm9/chgyYsG1ReSGUuW
YTySueNfWsXIl+sdb+lseZdqQWOuLcetqdIsoInHBlPxXvh6wCwwvDEkRNlNlrwH
U3k0mRuRTS7Ybl0PorGe+6Qm2t/wZnlZdH2B4NenBCcIxN62zcTd+KP5sIgi8zhu
YFMYpMY8/Is10YYhixK3deVPq9xAqYi6DvBX/aKrbF18Fu8zrM3nWDDGyuEUp6RJ
v1CuJwoloeQQClfN734DcXk3spJQONtwQAl5jn8bCCI75U/1N5DMrc4WPgaRRW+w
/ft4Ta1ReVoZyvZXlcURUwieVJ9Ldzvw9fTjWnoOjUAhZIHU16vnxLpBXf8HrpLo
tEd6JHkv0m2I/RqxwFqtfOX/ieGBtIE4FjypBaF2LgsNWfqciaEbvWX1XVLaq1cl
xLCqRhl1d4l59vIAlW51m62HKJnv0c+LcwXiJohXim5WNHnS+le7gJfzV3AUbIl9
t6mTjAmN75K4ErF1RMcqr5Ea8pO4UzTB8p0sASrmvdYEGitzc7fH2F5IiWMfdM67
0k6bnmYmhP4lA2U4uPHYBvo1ZPvIJRBA+pKwc33neVUcQNAgHLPluiTBPgNpZyYw
7c22IViKKuPY0F4DCB+kDqknzfg1i6GKEj0bb+7ydQHNhtOFmsReK1L4lF7tYJHx
4QATB/G7z0jKITku2cLyK/vzF+xpE+5hGlblLZb3mreJudmvOdmH+KN7A2gYEoRH
rgB3xkkQLH08pwr89CaNLS7W+d4XXsP0cHQ8sZtmfCbkMRUawxFLkGTSoO3/u0GQ
TfadFtT7ca0446dEMOkilEWH2rKqbmhKO6Q9x37pAxdaEcydBo8xwHmD9enHvG+w
zqi2k71EPxvcrfpa6fYKs6MKZgAarxUjKHYZvQS1hXO7Bm5vQlCB9zb7TwLaC7oM
RnTinRZduPsgtWx+ht9QYMK9z3grilK4eI31gc8M5Qz83idobtlP8s+6KdJD3UT1
mpmIgXK8o7i0o4cHdjBSoNWZNTBricb2u0nRis3vSI5Lw5YC4prjO9kQ8Zz7NYbO
2aOjTnNZppyXV8QjV6Uh6FXUCPpu7qYpB8ZwxfTOdEdhYCRu9yj9EIw9sJwjkb70
EKAy3U2yVAVShqlOfNcH3oWwZyqd1ITs/9RVvS+UyBK7AltrWSL1RnMyWMehrsK8
bQEz0fnromCDFBrepte6AlHYt1cVbGSw59KuEnubGwVZj35t9I5tLB7RpgCPg5eQ
LYySz84hndYf2Ta053QxZqw8E/6vYuUmgHg+qLCip7iGbQxl+8lYQsrPdyGGWOVx
JlKs+pGKG1MjhBM7Twto+MJvkacA9iZTK9AiH41Ppl+ktVOsYNx/eb7ZxcxMJlLu
TzYZv+TLygu7aB8eRcRovuLYfRcvNN6UAKO7N3l7KW/kYkeZ9O5y+NPVlpc0hwNv
7WehI7KIbB/e9/yNS3zuLg+iKTTs4kBXQ3O1CAyGJFkYrrnBob7F8KuowLVBS96z
dvwKaMm+YD+N4RB0zHTmF078Bfw5wKy2rLGev0piW8irjO+sLIcNh6ItRNgpHUIu
HzYMO0qjE95lr6cumaCLkomHZ+p5e3NAR7BKfqY2mmlbcWJ09qN45WDtnL9LGr+p
YLAR1GArA/EPB69rQPkRxyUjb0EqOvgjThxi29rRuQfA7zS+MUa/aiZ3yubl8qYp
3k0QBzD9PL8iPn6R59uDwu4z3tiZZqU1q668j1XVWGAhgIioLi9phZSu9SjMVnPy
vbVmWIDg5/nJ/LdMJIivsLFIVEM5fzxxRZBqv/K9rQrG8ULJHQT8WnUHzu3jiTSX
XDFCjDGBYnPOqoq+Vbn0/U/f+gt7IHm4DBIb+ky6qj3NitDBeJPZ0Zkb9E1bLhuL
WINzTfv6L7xfmXfsZdN+tgHWYtb7lsWxEr0sxBCMGwaesi/CRVuBOUHePeVtK2E9
t29oEGlHo4UOpLIQF9p8MA8HiAqgfrcIMjwnZwqCRnEKrrQWS5Uz/YALoWcKro6w
tQcNayz/14i4L77kN84y7lXauth8oR9V9v7tomWn0OEtZjdBZxQal9hepQdZKqTs
7XQnpb+XMX+fqrFFswenM2UTz45LzSC3RssAhCaEHxh3q/ymcNNLNGcognoesTsf
euFokO1FOYe2kpZNBJb7UMNTAy2CF4wfhkTAYyCB65R8ShO1+l1jKyYu1eOiHLS5
goOvEzdaGc5pEMTKYEML6Rq451MkdrnMMotok8vgqrdEDq3LSgx6ptKYB3ZjKRvM
FJxk3QQeGDWcL5KkP24ZTQsDyWuTghDTekkK643EFInscgxP7M+6MgCAuH3g7koR
HBEO5cJv9JFtB+M2n+3Y92TDWwSi/Cs6xN2cX6MwWEQoJ9axHYgEgM6rPhcqBnCd
1aK2XLbjRmjWN3X3f21JStBb6xkUh0ijFxpMXcXVnjuLqL4NuwwHpOKJrBviE45w
VDgn0EYx1MWMbx3x7tnCwHyUOiZPPHWCKGaaW0X30dZknZxODygpf56qZTiAf9su
Rs/y6zzsHh9/GMpyCLc6c6lX5O4V1Fy2RRFPnPX5RdhxYyE/LFg8ib63zYLaBKTD
Ds9cimfaLUGtLxd62bwpheNTpniEqSw3kVjSn4+NQ8NKWCFAhbGt+APn75G4WLMS
IF4wU4HHzqUVoPwjpiBEozTCyhk43inumeSe0L63jjdFKYB5+/zy+/5+c8r40ED2
iTRzXvR8f40/9fCa2Wb+KxNqfIu8GAQ3JS7UyyfThKkT+kVqwlraY2IInEESYVIc
XjeF/a/vL1/3vi/NU7XtEVxntRGrJowOFcjm4aQvwR7Hy77JbqrpowbJ3IUtvGlv
4PWsrWleh8BOxAYQV1bDUi3kD0elcD05OjPNOYfNwAj16lFladNRTjPKm2jT4uHx
8LeDFTqbjSL/+NaBTVU2XZ5UUsk5r3ERuPMer+fDS1WAYkckcbtcny7Lvj2+pfyQ
mSxqTujebNAtlrlo0R1ifjFVoZT12EkzqsuwktDCfHOFENcfEE0+FS5A4atynMHj
8r7lFFRPauJgCFS1rU7rz5bdG5lE8tY5Scfz4w4k23hIRcYPvnfXlmr2UrkjNe3c
edpIWvr0yHMHufFdDEk5avmATe4nUACexEAa3jGynXylnikza0EjgGS3zlw1XUi2
K1b8oYk+7eVoCPxU7wyLcaIdtehARX9vf9nonoO6UWgPiB9JO5P6mjPqDxqJVUak
xzKWKD4cAMSpAy3picx1df5eVBrR9jPqjqEgdmc+sP/hrJpjOxa487/lhsoCNvH5
p4/ChyNNczWe0IYU5/X23t76gmxD7hIcup4IqkjBiTXqxM6P16cDJLDMXYEhPZfg
iM9N/UufUtp9NrPsTXBCBtV0xZEyY7tDBCYlbprpNNTMu/I7Hhjp4uEteYrHBkUy
1LQi7x94S6Ue3Lhs/tHdpNrCOqhoHUMys856iKt9AZ5aQPGp0z7VerMy66Vo5P1y
ENvJvHvmv8zigr7V+RK+uwYcUZsY962q8jAZtAafL0INGNhUmvcHxIFZlefzTgui
23Z91eUUvyWqWr469W2piypyz//iP+TKS0ZyvzfbEcSA+Td9ytxVoXU8RDJC0up1
8IrzSPMl1cW1G+2Wdwvy9fLmH5Iybr3B/M/TlIf2/sC9QM+PmU8UoJocFiI5zOBE
UVkUOCwOUpVuZyW52eN0Q2y1hFIfbhL4O8jEFGQsjGm5FGZs5mIlwD/jTpSha5pW
XXyH0w5mE5uBKD+YfK1QvF88/NSVsv+nCI4ShYBBsPlOlrpJVwTgfLcD/SxC1/ck
ttlqmuCjqKmo8ZWD9qqS7meDcSKX1CjYfxTEKd9/WA0dgyT5b1skVspjQHzPf2Bp
N9wuQXz5Xg316vlxi9vjGeDAHGwJj45WhOAiV91cStRC+JipJRdAt2V6hWJToYNU
aACmaTaUB7mtgf2lm8ZFhUaNLaIaheOHd4sWaPF+caOoYQlVq+vVZ7VLnn8CnXw8
G94inL/J5ZUO6XWwRAhVBVWuoJy+/0kCVeu7CgMj3ETfi/k+xIamoLajdzh/6U6V
1Gn3q2bgs0m0Mo0rLNClXJMFVPxkl3IjL6Yfo6PNNObVHEDsIDPin3UiaDcaw4Sw
BVR1lQN/NWcJlgo4f5+WY75oHlrXJjESA71kev57sIKAswzVExoXu41vZNlw67cG
U2fJv8EH2xMjFlY7fl17iy0YmYo5jafVvzQXMnzzH7CXFh0tB3HRZO63F73H1MKo
EhCOXNK35ZhDtUjdCcbyAPGOSFmbnPEZmTHxoPbSoHHVaDgauuubRqDgpPBVHvxB
O/25bOkTWB/V3HZW727gWpHBmopux5XbaUKNF27sflthzboJ1hwp0hEN06L9epth
BxhS4tMZOKC9+COrJBnC65ekm6ASussC8H3uufkLcnA5Pd+IpFWS6Jf4AJXjNgFa
u0WMGQBRoHeen+VWfOTR5Mb610ao3hm9O6HmvNhUSXdtVANQIEykXjT7Zxe+oeg4
v4I95xHXxb5aIyeed9UA5ReNQ+qPg0MWFJXeQH9HU1qxb6w3okSyUYbxwqi2NS0J
WMwLN6Tzn/85PQYAcLolzXJUpCTW8WvaukpVXlgdLsQcHXhX2jpmtZnejkN2vv13
8Xm3uy9IV0Slj2ebIU3i98CUnw38A3F9WweDE6VVTYlYX3Gyayrh4B8Os3vanwHM
xwcRO4T1+TFMgzzbx2XfAWRFTZViIfxoXCkQO5+7uaTTyY1PEWw/INdPygriv8vt
NyYH48rMiTiS3BG2nTLT2X1BJHU98Fl5g8IlgQKwtncdzqjE+kiPCa+m4hYtFuuH
2l3OCDzW9kltsPF4Bb2bV3Yrx3hFlNu8YC3c223ncMFy8rpka2LYuqg6RIlEA6Oq
o9c+yGBm2kQrkgNxc/0PcN4dw/fESrp/TU+/uItY8tQzSR/7kgLyZXQ2lMDelQCS
CetewpWZBRFi2Ud1SSgVnJub5OtOXGSTc+8BPK+sQXph+iBIZhJJx69tzYmnVHRY
W9fb5PFNNwcUSglQ+66YTV6Q84iZVQdBcnpyCZlE2sbM86Sx1z1sQays/HgpLGi0
mC5HOQq6CgXU/Y7RTwKQztEhkf8p4F0adutO3YMDnydaJwr6WYhXjR8V0CnP+NZo
S6GuB9ZRDeVB/hENuQSsu8AcnoeX8DNFOw4bTeSTrkpSflcfJB7fnidq9jwhWNtI
NPd/mufPBOhuATtWriZ4VyXK8DycBjW2tBgdkBnxzOCAEJiJZ4I5jMK4yz3VG2EI
Bu/KYuEF7HvRfBOu3RQh8gn0sr4fYWbovDxVbO00jlFbVSSbI91WxbOXWKyHpAvY
FNIkeOLodMAjDfw3wwTPHNRRYewH2Wm9Czw+zaCvMQTu5wgqtyLdsPdKep5suvee
tnIcwdBHkF6LUHtNUHIOCkL75083dIczDdA9IY3pFAurnKbYd3EBPba9MSpbzGUL
1RWNNcYkLnl0Uo+w4KX2bCse2CjLG+E0gwa6IX1yIc0XVJntg/kjHIE7ziYykkNN
TLZSJpCD/72td9xoAoUpXdySRkb+EBZ5/Yr0FQzBA6wn9jN/HdULmZZvX2GVOY9D
TxH9ktqpELmC1gXyWrh8a7CoNo0oIueYnez/0qIp9uyJ3N9mlTFi1QX7v7TC0Tn4
K6GIBpQiMiwZRdzzSJoE0kCVKDmztXAlP0ZmURWlwUwBKdtvpvSTGhKkR8Wcgjka
JkpvFzlrXostLKBayOjxhagEmmzrGK0SQwF0UTQUUDRJgy1Ip7F4YrFP0c2LUtT0
s0nopNjDkFwGJwaOxhZVbQ/ofCbDO1ZAGiuuzTLaRl6z3T/8bZ6FvPGyC1STcW0D
4nSSiaKccR2ejNNOC1WcCjeFyp/d4sMFOEZcdE/IadyGAKxmy0SwX++jvrTzCSuD
6G/Y5BZkEIhuhFCX45iCTaSmzYJCDuHtQEDUJFs6EBZ/1N9VL/tA8t5PODN538g0
FZi+prK/5r8jz+WzXatBgOauOLYzxnEjztaV6ZHjC0m00VoFxjqTdAR0jZEijvIP
teohi/KlzpCDxCKidZWDfo8UnZk7tqm+p02DalIQfDGSRuhTBomlqdFLPKNSi8i2
aTQ5zqiqi9a7C7UvkANlgETkGsO6Yqd6sIVF7ALQW1EE3682ZFdq87QRQZbuuBFr
j8Mtlw6N0xDokBoArvGQTbSN0ZbavFHwcinFR4m9W+uyiFCBc4uppsJpa+Q7ZVXQ
m/Pv5CFKCsmnNF82IgjxFY6GeWb+ihT2QEVqeH1nkHfSKH6/JEZKwBskLRFtWgDI
HZl1kqZsgYL6CbzR1OPWrS1qabeL6zM3VRkNTvX2qoCAq5XLimgsBnkB+WsYNm/a
ejh2gtVdDGsj+/xfJ3505TK8vEVddt+iZGuAnA9euW/N+xlwq4aM+Lw0g71lsIAz
Vxv8lBKTS5XWapM0NPnYyB1BA8HqvuZNSNcYlYEvEyXDXNTEHEH4jYi2mB/OY//w
CzdxYe75HpTARZMf87rsM3MWGqpiur701TQeOsaPOegdjLwZu6sJAc29cFSrcD6Z
2XYidF+DP5QEyWLpk6zAgNJv0Al4aim17iRFc52DGR3tKMThueeH3p5KlauGCSO5
MDAm8FxB9LJB3sqR99q5CUAtv+iHNFYhIhdcksPCJpGiIwm4I8d/XnC7y40mZ1Lu
ju4VppmWBMFHQ/fhXa0cAJg3V1SplkmiqvlBhC7meuGev2BuJkN9yukT2pJbXlaE
ZE/hv3NMF3jIwnkR0XW2vZZCZj+sn8AnbBAv3f4bELIoykXu+2BWXLuf4TW7r9H/
4/KQwNZWy54tZ+8B0QE+pWAc8CePK1dNsKBj8qSoQo8vvTPqUja/GthkTP8gcGvA
92Cq9/wKb2Xa1RgqPXTyn7LvjJjcyuktaHJ30WxhTHoBSnNX+qm8iOqS2NWA1tCD
febm3dOAzneM5wHvBJw2cCSRfjoIbp5Fk0PzSedP1uH41ZOAhsSwx4m4iZUxPb0g
ASxt93l6UkWCbHahU2cWfy+QxuPNRFduHJh0+yxS2xF5XI3NYdksN2k0HoIBHKM5
8/M1JsBsskunBFmozPn0wGD0d8mF3I6HSAud657DiYYdXFmdQ+mHoXELvylt05w9
qzf4fEcN0emCZkBbWZBQ2OImvqcTK37IBEnA2T7OgJGn0cZWPvUel1dm0EmhWn3F
vcjZzNs2vKUnRiG4NLUGRb3nyv+VPAtRdM+lWGAOwz3+/PnjwAg7d0qnkBEuLAv4
ezkFRlHgtkGzK7KhjWJna5EoINh995QKZ4FaaEGr5uvIMhk/mB32fDGJGD8vv0jG
Br6E90uUJmOEa53CypbNwzkQrd4vYgLmmcjTQ4yczEsnCNlHBWtwSrrvWPVgo62A
QPZMrHiE/OKupyvwGtJ80dhrwbMcjL0gNEdda+emnr9XuQlLNVH05X22M/KwNWiJ
VnjKuZqSwXAhwhvXGiU07yq27G1IwoFozPcNkI7QWJvgKeHcgqKwQ1QoM8zflZNp
/2Pp33nv5HBZJtIrWVfr2Kqp4llMAzFKi/n40to5Ea80isKYzL3SYeEjy1qZDyRo
`pragma protect end_protected
