// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:54 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
QwmDh1VI/pI+N5YK9MRMd/gSGKaUj4atV4pz77VaECN+N12h3g6Jh+G7y/ifIVJr
QqKpl5GKu0+FPH/1QRXVdU6g4xPmB3cgSBXx2Pwpk6XVy5qFEZvNthzBSgfdFw9k
UCj73LrynJnSQ/gOc6AHXk86RaOF/uP3BhxEeZ+QvKc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7344)
/y0RVfEtq7WAiXGnUlCpsm5qNc/SYgoBQa+pEWEIYXwCtqOhfpOPBNx0yuIoWKLg
/5NrczZEtVRQvE+L/yrRsNJFqzRs8RKPomghUoLHlk89UbSwG2+xGZtgyVktbn/a
3bf8gWmTTlTgdqsfmBsGpSnkeYo+tVRPOlz8uSI1HXaVbJcLyHZJJCIKDrI83Teo
E0zI1oJ/SskoTmaNDg2JTnkM/nA0bu2kCU/4N2e5HJAqyi9R+TM2iF1mC3piL5M3
Rw308gc8QSJG4KK0BJlTA2P9ZZSo53irKiHu3JTEVE2wd33bqzosIOG35aoVsxrS
QK00JRt7zkbjAzT+7/LYu4MrHsVhh9q2mpQ/GTcfpGLTqk54pRQzih4WGpdagvck
TqaOdlFzgnEdS1ON4KAnzCyumjPekJoXOBey5ocTbQVrduTQcdahuvzaiOvowKT/
Dnb9Xcj4X4V08/HyJUa+bZC+4SanwpcDpsHZgZc/JurbJienCplEK1kH/qtRa6+L
Y4rWVwJu7QNZ/Bcltl49eucbo6IxIQFBV+6vhyFiCaF+eVoG2+GvRSpfgCsuEgx3
00cCmBdS4Y+aj/AirWseFVD1HlBBOF2B2OjWmevkjKqx42GTtOiotuWeJnrrLlTF
ZO6fsBCYcebOxqFOs/Ez26EQbKVFDRYZnLaO0sWymq5lXDsWE7LGTBa6SkH4DfQI
Y7feSZi6vd72bNFujYnGkt6sKNxE06RkvDE8gLgT949ImGuYoBM61+wGgxgCZ9Ry
v6g2qcYEVe2Prm275PUb+cInSxYHHYYRBcQ2yIlhbVHjo43TnEYH7eASAPWX5MUu
tzI6yOO9pyW/Zbh0L8ehqGctSDba2c3esiuOsIe1sO4+i5PR94Ypm0Gq5m6U39jc
0z6YxwWdXjT8HtKjkF/alhytEstzm3O3Mxb0i3mbWPgJL5vgsbedKivnpMSk7as+
TNzb98WJdocm6NT0yAS1oQuMwx5W7zgbwU/3+GIO94GDofF9gbHUndNV99K4Xl6K
Fd/r8T+JlbQgvt+ujUxbBQbKQ5pOuCyg2kN5S905Sfag9tBJMua3dUd92tzvxaYj
+SUWB0EApO1MerDiblPND24tIVk0iY8UecYmIMFDdzUjMWpR4yvP81ayfHmPxYsz
JtUR94mN5n7W/9mILCwZ3gKCY+o3k3B951W8UoimYhNywxCO2yDysp6A36chR0Vh
DrjWGH+MYWtmaXGUqJzjqJUhGCJ2b3OH2qRC4HJw+sW8v9dPDJCdj5qDiqX8rSBv
b8DVbiQZsSHOrt08GE0uEDfgtIX8NnIIamap+KSIbqEW6JAqbPN88q/PXqg2gOMx
/IzcfnteHvnHapJjLRVzxpWDwse0OcHRKmg5Rucm4woRBkpwfyAagQbaCWMKI0HR
dFLGawK4g0G6sP8HGGF4kaXZwURVZqbb2RPmwbapOkzMdRLg8DktdOOGMcjBN27/
xoZtplmqvC6ot5V8zyqxxjF/1DDr+xDkiBnOQuNKLcvRat/bYayWjXw7c89LeW28
uBRIBLcqlGqe+egHRsUw2kVanCycfSTQFSvEpVDa3DNpT6OgmIVWvMynsbrj/z8u
+zy689xcagkTXleqN8x1o4MauE1k9AXRsdv4P1Oku3TzQKiP/RwKC9fpzs5zFXd0
np7cCRYRRY2P6hYvGoNWWChrScACk0dB3UDDZr5OgFEVeUc95ncnSOtCTnt0sVpe
FP2E3OfCjgD8Hi61gabSdPeZTuJbuQA+oHhZohbQiu6x7yJFBkDCyB/+A7cTGgO6
nX6BcMn43qHdEsqpwuG1SkQ6dT+/jjkze8npBmZtSGhJZcrajexDuQqMSJwQBG43
cSaDXzbomO/4A/DdrBQxZmu0qKwykzhcyW1oYbfC5uh5Uaincw0aXEtvMpU+C4+s
KuSoSdiWeHEZ7O+A9a0FaryDMhFY6xl+lZaii77tKhkIdlyfNBi+N19D2i72XqZk
noDBxk7jeq8HrlVgeDgAPlgHjZ+Pp9VYyynXQgsN57BxchGrCVMMAn0DshSMgTe3
OOYZ4wa3tHVKkCCKM7CIdnCLJAzagXOW0DxSD7ot/0701RgBBCjejmkXmKKVFZyO
1FOAURQhGykp299zVSwJIFqe7q9VpTZkUAiWwCdreeWGc2TPzmp0fVaB+Bp//fdO
d8wONd7aZyplveBhO0T+IidESBSWn5Bq+lI6q1qZoMVYymgrx3a/uynNTZ2YlT7y
ei0zJAM13kphvlxq7MkrfuLkhKwP9l8XBqZKFJGWFVJhvFD7pQgo4E16wDg7ls9i
+PnLE3SypX+oDw027ddKdbD0QdIWTC8Q4Nsg8DwIoAQgARPREboLf/sI5DI2oFAx
s4PsaBMmM0S1/AfEoLqbpT/Rca1n6Vt9saZiKDWXyKizyKNqOiDOxq6BasdWXSwe
8ejt2AwmuJ4f9YGImHrkGkJKGqKAtOVObEQA1Ji/sQTjSbnNsr0xezXnfOSLw4Xj
gWukRPVwMR1MmN0brgbdXOm+KvkgGeD+io2PilU24QVm+JQv6cm4YN9j1xerjToQ
EP5bgPb7EqYQmhg7V5UUGp46t+aobyu9rdLoZZuFOWCbJI+lpBCtdRdAN/XOHWqH
ZLY0+J6KyMB/dM/3yRA3EP2dgu0VylXMzticBJlWNpeKY/mAEw9B7F5mYsksjvX4
axhGyVO/MS3gtmQNjvrCShlrHRgpuMbrApUDJ03Xd5d4Hefpt5aXpZddrF27S1P0
K6QioUoAC4e/hNB+1JE0447h/tZcfyyVeMqZZN7PLs7+H1RGrnm23qui7P1Vzxxd
t9JRIS7bNBRa3x9buBr7S4ibhygEw6DexL19JZJYCh2zknoKd3ns1UUzcjrqvtbF
MLDvxDfxO96dS8CSLJnkCC1MOCBnpjnUzitAuVAOBA2+x04j6m6zlPZu1YYDMT/1
1sMrRBN5vkp6a/gh1sCLc0KQaEdGq9VmBEreJS1+cbnJm0XafsKiMhYg4NmQe8SO
cwvqGlVRh3rL4tih6crthR38a8Oce2rxmUTwaKsbFTmQJKVd7TNhHTmHbaW9cX4o
fqs21FgTj8zS1POblALR457k/goEiyrGTfFCMVpZzlqUyVLGvSQZi/D1leWwZWOd
I2QFXbK3yDByP3BjMGs7PZ4DwGPSu1sQqJLhZT3uuM7cTCINTBU/b+uY1QEs95Lb
xQ4yq68c/jVbri8gDu2darXPuycKWtNjAVyQj4cHwMJz2AbzjO+ZkBN3pHWU9RDa
/ftSjtbqvK+dWoNO+hQoFCkf+pNqMCYVIu3u5ztdm8hCntUPgV9cDo3SNUYWRs9a
9tr2CzYQjD7QhbEGP3Rd7Rb6IVz7Qno/hovFfuxU5IKtFdP1xhb0CbxK/tyPcZ8Q
LXi8F8fIALI1FWl8V6NK5AbrGsl3FcySW50HzljCKGnD6PAcgH0VibaQRsmbhwls
8KRTNeudY6FdzV4ORhV2jB8riksiTZcuA65Ixhca9w0KPS8tJcz3cX+N85v11YM0
vvFCF88eSk8k9yl9HD3z5dbpJJVxx1+MTWfttVaPJEwiDcZoLB5tooshkoWBtAJF
hkQ5vOihcl3Z8/V+qyK57ZP//KUh6mdcPASU6prKMHXkoJJPHJ4u6/RzJezXTp2J
yYvjKPv4sjpSnLlEHiaedqJxFwslqS2NgXAfn/wTpAy0Xaf/uLupJcyvkXycorqg
t67TH9rDPuhTaPWBlumUvbjZq6Z7lfMN34oNJoCahQXoy+fJ2TZFJErXDuQRk7F0
e5CbxheizDy59FvpPCRLxtlvvIAQxqFj9DUAvxxHrPeWFFi2+8AX5VetCDeXKfqb
s7UAqjJOtmeTRIFIwC/ezKrwCigVkNjDDRh3aEGNdf/ky6hDH295FYDKkhk/WIyo
pP/xweeebqjhzVvJhI8fDLmXz88lAD1419ejCC4nnUWYXmeb01Gu3HigtVSwkS9G
HlJr4quLcr2OPAq+yVBIX6WQD3Mje6cZ78OsUO5X1MCV+KDih9osYumTCNn0IHM8
sYUzfwbLd8GEP7TYFnl5+4xGkJ7Eo8ghN27V2yed1Ee5KIAupKMo1EbQZU97HIv2
zXDkBgWo0q4idPRm9ujmUTloFQ2iVxLZPHgwiWjMyTdAGc/y9cg5VaT9PTfuQ+nG
GaouOGrGLQM4Fx4wNbWNGeZW1mCUo6aK+AQUJNLzkGmySZyqS/CHZrLQhit1iMK3
j4uCZGr9730Q28bEQHTY3WQSbG+IelByCZJpES6e+2vAnMr6FY9U1L5o6GjGkZaR
m3tl1jqkOf+8veOhY+iy2gJr6L+GzMDRgCOA0K+EkU+q7X2CZnZf5MRSWHGgj4bU
49ftNK4YzfW4+2lxWYjKiOPr0MdIMSXBSJQuWIKJ9AMzgpEyQs7Ow7rk52A1UfrK
0dC+zQHB6CVYODWn0FPbDA2mYOZ/eremKeR3HG1yEawF+d+cYQlzBVY3yjtWCDtx
eqVairZ6ZvPhxr5E0OqCneUCDeKXFCG9xHnFomZQK2bwc8D6zzPvk1bmq0gUpTnG
odZ/CFeOkXb0e8pJBPR+2FtwMu+yiDbxhhFl6gSkHMzSDUUGjI3eIKkwi2oLB/8P
MUIDiaON5XVx7Q2LrbTr0AIxfYNugpPG/a/kDcp0MvdafluJgGnvHrBdW4ml1nnq
7Acel5dl5xPTsWUhQ1for4tyjRhzxkWBRkhX8XB2EQ0vo8SPRFkpqvFW/q6Iky7x
TzKd2Qr9Fn6ubkICSJcmK0aaERHrM+P26uDqoXSzv/2KWFDKaBSvyv6jBBWKtRgZ
u6U4Ge6hEsvzsvGOOcZaguhT0S9cSC68X+N5KSoMzzYMV5KJc7VgB0h71VzwQ4kj
wJo3lbwyKbtaqoQFy/iPMgaD48EuwgJ15pgCJged+5rfZSom4Q89Z999zxTExiIY
19G+rlniU9C4R2Midam3ZsSwkEssL9KlX/ulTgZDxntl9O/14u6ESjoZe8ccnfzE
DlD4oNxHrxDUvjI7zI1vX0q4+Ht3blP58+QdALYg/1+XsDypy/WNRkAPN7/wNodo
mNWrW+6ozo216d6RzpWlBWh2DQdPvBswEmMgjIGkzqvFf1GBpS33boO2VnCaDkmW
n0wPPUG+9B8wIZZqGLs5f0RF7YZjbmdltuu0PMv6lYjj/W3GMb6tRSrLMumEbDCq
m8qNOqFBJWeK5QssY5rxfeoZ/KExJ2KtyygjxncJHkWfQKaGKsKs4LYD9juxK/9j
zF8Qb8isU8TkFkbma0hVHQL3b9q6qtsFTEGmCBnjBSfku6fHYTRxN94yJY02qYeN
8+XpKkEyPlfVkmQDCYCyUckCA2SSR+QaW56PuZVI0ic3bsqqKNNaywH1jkCVnNX2
1Ms3RAhZSzDpIFqvW3iLTpDSKH/+g9meJNK1WbBw7R56o8vms1/QpXN8rTf+kdVL
am3iVlBfvt6UQKLDC4g/aab+g4IWYXTEJUbC4ds+yXzTm0tuMavMtRuOhFNsJ9dV
4ijUzL0k4/ItbLgLpwF6o7HbVcj5r28D74e9EASnEt1d1/7BGlthnz7XeB2JigyB
Q/jR672BYkNFmr+1lkt96RV1+FliICHDqeupOMcz7gEMNNWDmjGcyvdGvvlzAga7
zprkWZik16Jeijn+JmY3VKSgjhiDw4TX4KUwxtYsDmJQu3bzy78MBErWJO4BQeHE
fh6/1RC9VLg8sF6ozLD+BEak8UHc0gkseruhYAUvH/nThGwMczcaRhuMvTTLsiYq
LVnHsLytSSQ0Ekn16m96i+tUBChJetuGTgd2v/7iPvWHxqq/jvKIav5JsgFMth3v
NLKKnWWZ1XoPNAitOh3htjFZxyiLuvTzITyRAYBtbOGXa6nO3MG9f6BxPiianbWd
YxX+yjM8XohBZc4hEA7sgEfrU6/Ek4FqxzKrpibhl3X0BLl+21alpcsW4Vekomta
rtqTKwUn/GbtELGqVkMgBG/lUSJqh/CxVM6s94XLVxPeEs9M/3rIrKElckuQthkv
8nnpJL4wLXaRrDpFblFKiZlcAVmr1wDhAssTy0/VJ8/W/YuTxaM+eHkPAKIpUcLA
K1NsI1feiIzhQD5LVHcJqN5Cq74DKCfdsjMlKsZypv1GiZ06JF8wdQ1JxbwLKEGB
mI8BL31fvWmxftq03mdStKOvLSJH8Kjq6jaYOzY+MgDRue7wUeDZhbYm2bk1h0RS
1hWvepbJSmIpa2L633IdDD7/JUYaBHqkC/Jox5pMNQ7Xshmub0yzTqKOm9V0UttF
m6c0bAEIs+/duSQDdoJ4mm3Ok52B0QWnZOvXvL6f4yFhfRxgnM8260e4za8jbuip
AaDKpOPDJ09EvQyhJ/+wNB7BFTHkF4h+7QWqfFkr6eJbdIXYr0esCjMJlfB9JOM+
aEBLn6CddZJMbeLmq0JzZuCC89UmhtWVbL+e4xrfktbeXX7C5QPhFJwyvjTTbn9Y
5pnrOzr4ZYxwW8kVAqQJRwPgkdAlxlM/jLS0OvFMZHXalAzt66rapleJHBJ+WKu6
Pin2Yj1CUXrayBoEhSw5DyLZ8Oebqm2OEfi9mR/QLDtsmDPgEpW62FKlxmW7aCh1
96Lq0bPR1NzAtMPdqPojPzgvpw1RSjiQdisgQsR6uW5w8grZTT2hwkNAsiX3MQpF
e6dX8bChlVfXBPxGiEeLUmqqFsoEaj+TYsdUmE4y6o5L8WeDJl7ABVfCNMbbi4Zg
lg8WZepGnZoK1CEBKVU5BHnhRvuVfzuQoy4RiyDk/plpDuved5V+swIZOsdbDyGg
AmFhSz/0F4aCNniALljWCk0O7OikBrWX/fYlJI1zY7ObfxMdXxXhNjlxMhs7Zmj8
90U4DduLZZyMWnSE41LnZ0sIPHueLATu2ly/SP7YNjRzavZwC1/0Dtm6y0OPnBdZ
QwZS3p6MB30Q6Vcmot2LxKnKhloyZIPcUgyAl5RKBdYiF8nUGtiQq9jIm3a7iJPP
/t9NPQ54PX4k/fQFJoLc1RY6E0PSikwFWQn+mjXmV72nDtUvEhU6XYFwB8+6rWk/
iicylROuEwJpcHJYGabVM99GG/bdkF3lFyzi4TYHJygaNLbR70GLJmfHKyzVcEWZ
hIqqiKFXsilrEZApbI9l6rGYN/My78oRpfuMyqVyzuAR9JfkFYlCq18OQIDSE3J4
VztF6YOC/nWGkt49s1tmVi6DVcgLd1kwb/cWqvxqBByQBcZ8uowFzpWXYpTqmm3E
aa/GaWRnx7n5QPFR4POwHekrGER+anFSv3BUNOKxVe1GuwbaASPi7Wc0kR9Vu3D5
wz5NJsJuvvQ3fn0q3+LyXC5fKgvMXNv538Dgl9oMkaUxP7XShHBGc7v7+ynSEvdv
+Mt37V9FNTcEHTwcScLxXNQd1nti7WkqEQxQaf6MosuDZvPMRVinHMpalmeclI6Z
l4ujvDxd1whwvG8vA6PuPbjwrjzD8SFhRl2iyS0sru8mS5Od+llPNqYmhnNSk97i
4tFCrE9biNNrAvS4hEwAsGazsb55Q0Tvo+RIJIP/I5dhMunMd4vTqunkL6GOKi0/
hqo8pycOO9Q6AVjAiWnCy19AAaoBnyBT6VygPChRtfjxksA1BAd+I9TiYIcvqBN1
qGU2PWAcspA8rG73jJe8FOU7NCuc41VbljwEPEDMoL2lj7wVwTNRmrBzgeGm9uGa
mJiqB0hgLeVWS5rTigJ76zRcg8EbwfP+zsjj0pMKPaQftjKILZyDFPAnIaCmWG5Y
QdGhrCM/WybzF7L1hu6VqeMUVD42hWRdZyMHR88MfoAhAoRJwEIsL/PkmnV5+zLr
zOfsKrfTrYO+OXKBcJpX7Y/bXnBZsnq42iyEPPtqIXBGUesMz/zOIYVuxun4Em0u
2EJuIAWudQAWfioL3u6s9y6OuUgTazUnbZqw8LlzTeS9/hpW8TevuiDHwl5bS1n5
Z7L9lVQU0LxK3wEgQnEqjcYZjADQ5Fl0H9ci4PUcJqbe9kyqegwQ5S11d6iBFXG2
9TpeAbDFFfv8VN4EPtYbNwcaBkKAesntK1iM6aGlVtSSxMPLeowJTvgqfWxJrwAQ
RCHuyQ2aGWuplKmRnIS2l9vrBDORdyRpggZTWJSPTujAwA+EBI+yERXbCOL8p9A7
zc/SlNFempN8OxXUyp9MuXSvemI75q+4/3vHnNOamo3ZmnOsveI/MJPyPFd67lNP
+u+n812arA7AGYyfhCruj61Fmu4cIKOQKfWnR4DbwnEZooBh/aFVbGS2EZMoPOuh
ziJf8YRv73rT2WG/h8txDKO9yKD17pUuK/lJ955n3W5IwGTommrDrkQ1G/4isCro
0F/7p5JCDeoZQcP4Bbg10ZUxGBIFHBW28pQ1HCueC60E6ukVLeCiwJI2w7SCmNya
nFFpJ9TeAWOdYoKiddXd7FeYqnUz0WwTsFw7drzfl9HmWGsD8WtPV3yv+bSpGzH+
+An17lspThGb88Ao7qOn9DNZ2/ZvinCDXc2/1iDIzFohIooi120KYbMw9YWcdosS
3MdMndvJlyJrcBEUMD5pP3XZ+9BocAgNEDwhF0idmc8IJmdXlNAkWD/Hp7tQUG/C
H2VeWYtLZ+f1D2l59c8Fm2oN1L2vPtNbHgj77UDScGwr9MXwHMR6hd/lHBmPnPIK
vA3lsTrzng+c5RIHJveHzhsaFKsKSibfJyaXEHW+OUYCAity1ufEWqcCIH/nnPWK
z35DbduwRtgF6+d/3M5Zh9egnE1PVeRKkpjf6RNsn141quVMOP+GHh1fhi0Wf6pO
N1pwpegzerwgA+/ToEHWrp1d/7f4QsdbFdE/1aDM8l1hOTViRKBO2mYcD1zkQLdT
BWsUy7EvG3tmKAzxeaZ4t2chhNEP/L/FmmvJPGTyDxLDX/6IDjPkz0Umf3jW08g2
FYboSb6RQ2RjdRJ61J4y+AOZMJ2G+zmv1C6nU6UpLdHfhEA/z9HctmA7of7aGufC
I9Bblq8Mwj/drGC7iblbbEG2Xfo8fWSIEwXcXaLWHTo4XOF3WJCAJ2It94GhXyqL
PPrBUUZLLgwuanEzzrT6LKh6rJ+HivaZX1V4iej5hZyKx7K1SV5bhuYLZvwGwhZ+
JcJHCxTR5sTFBsoqHQbnbZRWx0v8GJ4lPUgwyMDz+yHkcs88E2xz/M4oSHtVu049
9OCQa0hSniG3GnIc0JaWBX3DQlwCBdOGtuwyrhGpsd3CNFzf7WliRHkjUe0UkjLZ
m7IMai8JkdMkzEuu2YvtlbVUQsVY0p58rk73fzbFIMrt0Tyibh2yZqgQct5c2vlZ
R+pWyIW8VN7H03X6DEqhiT9jnp3ivOM2PQlJj9U2lkqaWdk5GmJ5QVglc2Bh2TrD
RXUSzgrwqqSU3LwULUNNGTtjRcqTYsku1Fjfwv53DCsPaRb3kJXo3dmvuPq6XSLZ
CLYJZ+O4kP8TsDw+6T5S8uqmAH4mAwPhvWHwLB9tg7C7T0iVh3grdYn104UpsxFH
LleexoFAi//slkU7YwpdcqxSHvRL2dtU4ZhZG50/1Mx7dRRasvcMR1jwK9PdA7jp
HE8IfwOTpA/G7A1vBCUGS7AbEtqpthrZyFWTwGT4F0ya4fmdssqmh4UQ4HabUjZK
QU1goddogeuDL4bT+MkzUKFyeYsoFiISZmzkoHGB/Lw9pyGFbTUsO8zkVSrHgUZ/
8jusiCT7ihdGVDHPr1Kyun91GOIpfO6EqkmDJZPR1gsqGUXE8A0Gunm7+Na8zABN
2MMLlNu7OECfvnB7RIGrTMfxUgVCcrqUI5KW/jeTP8L1jvnwfnBqqjxQK7CCVyFK
`pragma protect end_protected
