// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:50 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
qmN9oUM5Y6ARKMRv0xadw6nZR9a4NDGxUpUrm1v9WQIN5/o1Se8l2W41QM70Wkjs
g8RqGrTaqz2U0BWZrQsl2VmcwcT8vguPs+VTXxAvjmOclCOLDe3Pwd6uZ6UHe+PD
/uEn7kcstZHYUaqEoFM/KJ2lIl11QQyO1MKbN3mYrcY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 82848)
GghvK22XbMyla9+WyHhh+HHCAQm9B+6ry2BLhZXTx0no4pEglqZAGeGlds1kYbNb
rPjVLIbhiXgojO96NCvE0wJyXgsWJzBX3ZKr4R/b18jo7j+nwuEP81EXK4y2i60T
zYX38XiZmqrrcVVUvk+CSfbl0UmjgGrbj4S+kyPMCIXskCXGjVCTeCIBovDGjT4B
0OXQkibKCAYngRgOgqzNX/Vnb2+HYym1Kul1dVu05sLeR85boI5qSNOnZc+ZtK1F
/2Y2lCzm2dV2vyjNgzvIBlJMO1OS+oF/Jjf9N1Wwt5fz8G+rvVCW8gKjrqKoefV5
QZQhqJ7CbYJ/3DA1AbuMMA2C2K/y9IlxqerX7B9mJcLAsZFCX+w/VFyHQ/D43vSb
gffmwh4bYOc5oghO/oSxeXRZBDiamKzc05sSfDmyaAzMCWgC2BAMDpEGKrRtN2Bb
CENbuUTwHWqnC1DheinH3G9Ix04EWeK0laoyn/jiJsHDWnzMhpoNTav3k1cbkx4M
D8PDF4y908AOYBcb4s2YbUQ0kUUK5PhEyBAW/Gg8cz4U0qVMoqAYsIH84lzWYNwr
keSXazm9kFnibohaFth+N+YQmrrCMVsyhV1ZAXQYYzUqfHzuKLI+heIJRMZLIrNu
orZmqoWfszOZVwXrQTH5KBgplQ3jhaBO9M2lWleBPB2E16tycA4lR777JyZbsM8c
aAK8QDM2FzB4guW+ZLqTMgROoilRezV3ZyIsDlKLXwPYcbc6e6MFeEJw38uDbz/2
GH3ImDk3DuvJJAo1Wt9ZmOguDRqgXX/WkAON1wNQJEmE3T2i5cbtcAJr7bjZpdHa
SaoGNLbBEYvPDml+h+GSC4VOyOxImX7++C/iRewCL5Onw2GNcDIQkEMYL8WIosil
NOYzXfeWSI06YkPG55RuJNSkqaWflCsr7JcTjGbPHv6OecSCMYsknsMEsKqkLnEg
7T4KXpDsZ7K3dWVlonRAFgFmq0WIZ9UWhn50YtdImrpu+ahtX8JhtfN4otr655lE
xumK8xgQQkd6S2jETv2Q8nHdEgFhFGTeF3iYhK9gx2GvvQJpkYTi8D3Ekp/ln6oY
1e5f6Ppx2m9uboqZsS3zWSqlhnwNBQSRsbcZwP4NJmCG9jzs4AvmbEHL0V+ZixS5
WXfkF50jycp2O4TA7pTUIHnHpf7WboaP1OnHxW+NEHPpZmR6X6iytUmPnZE74KMa
ZkLWhe7ZGgQPpTtsEcA69nr/eTpk69FrjonRoRSxC0RshRT9yTGk2Tof40Hommpq
GK4K+u3TUxnuJuy5f/1UBUHOMmLdDv1qRYNrT7avOfTQ1cL4JJi6+Z8uz8SM3pdU
Etj6AGJA1ESoTdzmY7F+w81vIMbc6HO+gPT7FSAtwPQ0C/JtcTbmEMRIgIkMCCK8
ffGR3c8VZ63xT0xdCFXpsDWE4Qg1UHkStPXYWH7vrPhsQsBg6OtRh77Aw45F9SZi
YLEEiZcZJMI4pRAzDptjk8ug/3dEg73Y3b4nNVJDWPDmnZ/hZiNoTXOlkaGJ0Err
Ie8KspIJH3biVfSPvmc6xbxZFyFHElIjEspSbwR0kfgcC0CqqT3i9SmxgELzFEkz
p0XikVCNzdNyU84QqnhPc5glB8ampKImsHo/DUaApWoIVdTVYeO4sThkb/msJ7NJ
cki66+d8dngmKMmk5A0dUM0vg4raBJB74ltuzdQw5w6I6re9l+2C/hreCL1d+GSw
jK8q/q+3nk28b9gcDWxi7UVg6FuME8TSx21gm/rAhTJ6WTJERwGUPzx0wqhS7+bk
BWw85CWZ7aYVfaAEAVx5RqsP9fkGP09v3GQN2VPXUcvuJ9l0/ICTMGrU8vR7EiIO
xdM1Rh6MtysZ3c6MTP6JRQmxbPbGxhO1K9bVPjXosDIZ7iflfrQZn3uRLk0aC0VO
PxWFgP2e52WEaLVnt5S/PjvmHnSeCADDTus9FDMDJZqKqNdMPLll0D4j58JxImZD
Fct8jWbvAFAOEVJiIJZejstJ4hk2ALbKEAhOX8yWdx6URECE9kPvaTQo6qWua4fg
Phnjk4UifFeeLCZIy5weGCNeiO1DX1n1JBOjGuoK0F+gjp5wWVTT6c+GHMXT7NzN
V9EpEtqmcjTJNXnBXP2EZbyQtnVZ7jWCxOk0CGo5asq4ZH3TvY4Y6lpgYQyUMdiQ
Vlo5afymOiNq1aQChoxVuNicAxGO01F2xT85pZXr+5mYefiSIF6Q7CoBu0CYlrpQ
Sykajfhak64pJzDwk3shce9+gRC0hT66UPz+YK5VmJEiH7kfTxtKhnEYW9AXTIOr
QCl1M6+Z7HXZLji3CiTG8aA1MA5NuVx3wQskmofvXMKdDpJgHpbvBgXG1bvEqdP+
K51w4xI9lUi776+aJxsoSGInsbnY17+UlcFQTIs4twkmExi3TcLpKYy8fH8/p4cZ
DQuXkk/7L1MxOt9qmkhMX10bOg7ec830/CHkIcWPkbsu5f/VxMTzL5kCJQ3FVvq4
tinH3Bdt/qP5J/yrcWdbhxfiKJL6YIVddqiIBAalVCEtWY6RBSHTCeBLYbpjb+D8
BjI9QviUrayTGsgaOr7eDHJW7o+mJxE9JsdF+bh5QmO/0dpUV9mZPsP7g+aZ8Jmm
+sj1zEgO6U7ex68SnkAJWDxQUgr27CtOmXqpsKdf5gkfUBG4//Ycp6PTGYFE/3wk
c/JwxTgivYOl5VIyOvAXhr5lFDpaxqJIyw/eb3fO1LQd945rFx5D0xWEixiZPBac
WQVEd4w8k09X2zu0e4o3KLYQmVnlucguvPg2vcia2n6ai2ncvsDyI8BmkUyFxKTz
f1/o1l1S758pRVSiobVSWB39Jo+2Dj/zj1DwNKqclM1XUBGzt1eq8hBolFeG+SK3
OzW1V8hIp7E606NvJ0RAHN+Lx8DTTKeJNmu1fU5ytbeJdkXj3ylh/KIVBIRIS/XC
fEw3m80SnEHHI7MgF99iuIzzQSuLe9k/sl0SnvwwhMdg6ucq7wERq27YMfAO0qy9
ZFNQEET6qw0PONw1chplU/+2ke2h3hlrZJeSN0wrLFkPz9gUOi9dWSVe/ppBzRpF
7mbzkf7+rWSCUQk4zM+JzJWuR1NbJRrEtmiseBeFwGDSsi2m8zA0AWxcHjmR2qfB
Q8NJKLq+34iCiWwjQO7Ee7cvXh5jjXzIPnvnkdxhWE7rInnNKgOKRklPDnkK7Zrc
i3vT5aFfELYuV+c0QnG8p8qtfZ7oeXwICkxqjksawM/KnbfrhV4Pb7AWQBrhdYv5
ex5riOBJn0q7JKAf2yPl4VrqXmtM77vH4MJRfys6dc0X4A2es6ZL2LUVHO8bImSt
+dQ/qtRLtzmen3Ykerbt0QALhpZzJAFjWbMFfLUXkZrXqOGSyyJC2w1Fjv3xPqXS
9OHhOwNGV/765Lc8feYmmrj7uT7I3vmrAEznGgQ8nmmPp+TepJK4hv7QwaqSXayW
LW1Hs/4zlvegl4+arFqHXC/4gfMDbGgk8KbEW2onSUHA6k51dnyFf09BCNK5KjJv
AWGh+0TEMiJGzG0wMHgc8Gpc4jxV7gPPLOjv7KV8b7SVrVMOpH3FLGyPsjc/wdPA
WIbh7tRSZvhyLxciD5FMB5j1S5/OkGRe5V2KoabNrkDsr1Em8EkMncwFW186njoI
O7JgMIC8pnJB0ox5Zr5sqqIP/RZYmphyvEqzqPlrq1VTgMJR4rDo50MGeM411+l3
4D47xGVH3uRu0eGb5OjmhhJCXLTSnc0NdM7ciSfkmcFC7TEPZdEtSmW+LgJ8zF1J
j6+w7zhm29cfyfdVHChN+v1sPpQPHgrpLI8GYg0onjdmxRPHGjBl8/EDSdOgHO2P
L8EWpPf8KQHtMC0ZZazK6jgHwmWc/7uqQpT1WkGI9S5GQgZ/TzQrIBjo/eN1PC+T
rl9OPa7VYz9qbo8tXWljpwtQtzWr4kI1B5eSTFj66FPEpYmGLFQofdovROV4MjMI
K0d3WxvEfqwMoS/fhzRcO1rhyeXveVIl2Zrx++LOdL36bdMkZtLxzm4bndvCHAbR
C5soWJLuU1kyGVrog4AvqlibFxY16NXh5N6+6R3IUWtrlRl9yaLYfXwQmA+9G4fm
aqOWflmQaVCa85RioinxPVVlsI+XU5T0EfhE7skgYqhcDSRL3FuOBZ64MrGp9Et5
isDwjlg1x6Q1/X6LxCJj8ryAWB0S+5ugGzeEWve24SmVvnFZLbNae8XxcD21cbHH
5wb71bXgQ8zggd0PzeCpMh5tfhlOz3uWtG3dPQaPp3oj5Ser65ZsqEnqxSv4BHJ+
NoxL1WmRYDMDuXQFVsT829b4atDqIAQFPql5ssE2drvCtfiMbW7e5knmHBF7XJBk
PdESGL5FdsAc2IsLTjnFo+nocO7aXX3+Bq3wRS9R+3y16d6dZX6MKqXsThchskIy
bhi6grMJtLEQKrN2X2NpbJcvWq4IcLYBqJPZBM2CsnkJfN7oMxr/LLLPzMpm3ZZC
u2+VQfcKykCKSPTQoBCEU8SqP1rc99OOU9DtINddRzDSMaUKKeu9Y1BzxW6lXfPG
btPdO8eAMudhrC2tFRWtDtcduFZDTJFCAMtN1pF4E3I4OayYwI/dcnk5URTcgv7a
Iwadc53vS0vWbwrVYJvF3+Roj2vQ+FNboA1Qk7oIL985shMWZ0erUbvvhxi0FxjA
fi1+Biy3IkzurQPTnKFgMQaCW4tfrYWd2x3zewV8pnVq9uI/W+STC7hOMwvkHTg/
SlbAAg8LDbX/qHrWtjcWF3EN13Jwc3jUIgRonwi7lgpMBOnps6Cbxy6KafMs+sOl
A/+Ffza/o2FFTCIT/BOhrWMnJxlS+n9ZnU/lArjPwMzowzoSw6P/aGwoB6gGN4aL
jKDLwwooEpsVHF1XvWOGzQT2vusQyPO+bv+DnQy+MyUiolEqKDxrduISCMrzQ9Vy
SKph/K6qNjLcYXSipJRbsMI0Gj7nWk2vf4NwF+IJuyo1uRMhqW468QJxXZQmoZ2d
8OwLiFGhEzNkXoeQL56VB7yizYr1ynDlXbwXbokh+cPhdmrYyn/3rdRs2jaxa0eW
eGLgcmqSE1sETz6Iv/FPBt4PwuKJTvIUc1aTpZRG/lmvqSo2sBIMH4r6bhOcWK+S
J2KQe99mMj2a2e+q6J47DVmzTqsnpphCepHs7jkm2BkkILeLX8EIAyXZlT0gxes0
UAiaeL79Jlv6/aJusLKQWSlQlUDPkJSQd4y+ycUpheDDFWm/UWbHColOXQ25rLjL
sW0XVRZXvDhKVI45zZbOHUUslHQlH/sFfsJTzrSR6z8v45OXsrry9Lg+j8JNhVNf
vd3vd0giwkvpQ+o8ory2/UcYmIVaFs7j3zJuOnLSHTdUS1lZWBfZ38+BmPJRJmTA
0YmfPkQZ+f+rQG5JR6z4Nka/51HngMM4iYcvHB0GNTDXSOUjnmB5CCxq+AcBZoaB
vxSgV+iNCXuZl3jYIlwzOVA+5Ku6mx2YsT+63LQYmaG513nMz0Ljwb1dpblgx2Oi
VbjZVZeXP6faeeHHJcwmxmpOnG7KH5GD6T5uY1Iv07R9bLKhxJQmu80zNzb95T5h
ZbkguvkeA3XRXnyp3UFHtE4L3PyTnFHi+tHXsWwnRYzO+NfFGTZKjn8nuFCooJB6
4ob8Lk/ut0DJCbXDIrxPuYdOObhSuZ3YJauxZu0oSXNZ8BqkybEKSCL5EvE/sC0Q
Er3JlPoCXdpYKczAW3r3ST8e4JMKj+KEW3RYg+m7V9FEJp/kLOPlV9ob6KtNaGZK
goZWB0V+XNkrf/6i83xE9IRCRlOt8/Va2GtoU0htC5tOU62E6uE8sLjyt8evjC6H
X7joP2gwSaYlvNxkY/ZD6SGnikTr+xo9NyaAYMRPHhRWf6id5Ci5iT0dLv7GOwux
C9rgleWRMpkSttmjxXUN9x/acDIjG2tLO0LJWCrqFEFZg6dsZPOEENP44Ipimg75
LEDl7vJyoiXGJ0T6LHVwr+y1KiasP6HquFgfYNpuHmzvZleyv8DV5rNm8V3awB15
jfjlK0NqqoDYEKlwvdr+w8dEXgWsyGPqAwTFLAJ+1tyRZmYjkFMWVyUI5YL08hId
aT2UydyYJiOYLX0tBBYmV25RZI5uYvRxjmgihE15rh0O17bT7Le8QKwMQUmyv0aF
cUqpH1mKT6uh/2qdOUA02G3/9TUVTUx7HYNQo1Opn3hFRumDH3b+KkhT0pEL5rg7
jqL+0Jve7SwpRZKAwCClP7dg4kkKZV2VyV8yEA+XhQYcFp4NQ4w42NSxRHz8Sy5X
lIUdZ3Ta5NKLcBLORQ1zPJpLfLYBFIVvIkblwwp3o1Hv1vKr6HcNTd9Ge48Dy1Od
i7bJj0sEPQTzy4b5HbB8BCon5QXXQqk9Xpp1MQyPb3tvoJDT9i2kDCBg6MHMzdKJ
hmECkSQC7CwfzDOZw74sVR6Y7HWtWoy81y91airUR7xsK4a8xLvkeCN3XN08DrgC
jQFdehm0hxEaBNa0O1a0R9DWvZJV0ppJmEuiRLTQE/39p9Bc2qErq2MaFobNjiEt
S9Iq46v5CQpyTMCbtg7kNu+cx26ZAXF8ciginFAAHcyXQp3ZS7/XgBy3zNJHCSEG
z7xqZEaHfU0WQcU+/ulS57At2VtzCwXlMZkXQ6M89DTg2YRBrj5eE0P3s4HBe7h3
8U4HC0bdAE1fubsA5x52LZ/o07VCtzADzZaoE8zrEAio7QzKpyohSuXR0C2JFBtD
xsJGlmZY8KEtk+c0kXh+K3lCmV4ZBilfenKf2mQa6waY68wZbu17Y+jgVkONuKbI
/ycksQo3VM7jXOo3wAlPBPg84n33Ie2HN/aJsHd5qS8N/Hr79S1d0z2Vn+SRy27A
bY9CD/zKB1v1HOQCZ+Usx95d9mY4dx2tkEZoxR2ShBvBOwAuk7uZX4uFaJbS16Vg
z5183c3aQDvXthDuqRT4n1HOFxDFFGYcvgtso39H/0iTWNqN86DinuSc3Q2aqgYv
mrn1T3MW5MofGR93Kow/dhaxtZNhUqjnhbvX/6W7XNoPQ7xGqt5CESDwHl4oK1WJ
BRWMPKnKvdGe30+EWyX4PzQLIf00rRhF+qmf4jqc9TqAgIQFAZ0ilNBzopKvYnmp
aPDCF3i47TV8v0zXvYcnVogRnlVVeYq191nCM6Znm0SCCMpWwHoIW6l4K3Jwzr55
j8LhkzQ0scT96AI5bjQmgB2nBG2CIk1QGE8H4p8kxxnvsjul8UaDcUNJqXrOIZq5
6YQMh8BQXHxI8x3x9eR+vF74k5IVGMGY2KRrfEt4SndWQ8VkrbkRHR/ri93VdoQE
t3eX24irimw90NJ9qeIslgI6i0/EvNwmRurjHd60ybetwuSDN3MntqxxqHMonjVa
uey6lGldEPSc6TTh72DB8VmRdhMBFdLoKueEpY3m+m+iBkMrse6sx81LSdXa4wmM
/OztONUORC0vRqkNhpS7qALiwSwTRM4r9X8Au6XQoOGrLVh2pZMz6y0RajusZKB+
9nGjw9tlfi6eKSPuC6phJaqH6B/lyusH5Ue3qjHyo3WFfHD/TE5Qx3OaL2gTnQfJ
eZwcO8pXJqS1iYB8eBv28KTn04Dh10J9Z3rM5Kr05bCcJix9ji9aCiZokMm76H1t
UO6+ZfUcYZ4UrlFwCQOuZjWzq5diCREJoWqfAfiBsOQgPWfAcbHgtAsa6+8BEbTj
2cmjHEqD9KdVGoPrT/koe+M2fvvCOHIZVJycx6sITAFQyWx0aTpgrOE9LniXKA3b
ZC648zapBIB+C+PM5+voe3z1BNW8t27KhTzNZep6s34ya48n9vHVwjRYSNiDGCj5
zV1pWnKBfXUSQpeFTG30tkrnCD8BEipThOBSsvByPlLpH9cIRXQ6a7TfWy9ULlUK
gOAE2w8qBzgBFR+OOW1qpGww+C4pCV7Q/8fg6o9aCMYxeYNyMk7JEC38ou4cswy2
DqHTFwycWz9T6XJprea+vaK2pzbWLvuZ8/BBXKCsSFZ1ZsonVEAJlwcLtf66QAv9
azuFo9mXpyh0qgqvxHLh7G70x3cSFrYgChQNFvLr3qTRKnLla/hKchcJJOS0COVh
MU/qOGlsNAc5D/0DXqLYKc+ZtJMIOq5sATwq67h6IlRZE3IrsHdCWbfcMbRTOeD+
EHMPn+PZkaGPzfjd4FJONDxakTOp3p8et2guS4J8mN+WiBIzehzxRxFVoW4is65j
flV1pHCww/+uKyxzHtm1tqrA4J95W9AhF/mfceiWPudI2uGCgAbHYob060z3FOiw
OkdOhd1Wkv20V4ht8bIQ6rcOUBoew36pWonPcXHbHu7GBvGsgYOdwsmzm+wocHdR
kOGOtJfbMY4rEIyqufpE8ArmeWSevz4rKcEl6mz2xd5ekk4XxJ+zen49rKEu+tFu
Gf8FCttQWNe4O2seb2sEBLyWv4damhwpgpDXGvz/ip/SUeP08fB5J56jRrhTaQM/
XfFu0ouFUdkL1ZiUsHrQGFmVXGlTm15Cyy0pVIG0gbh0wd5xMuHcXvjO/8459bqG
+rYWPVMOM/dsRNOXB7uL4XUypU5+NwnMO9maI9SoHGWOsL6xcSe49LBE9325ETyD
wCKu2Mbn+gr6tAGypQ5MeLM8dMWez9fzpJLZ/fzRWOBgoCxrmkepn4ecYlGoD2pz
8aApCpU0nKJjg9EMVJKl7pft0xJ/UwX0Ud3XykajVhfHdNDL2kxyPKaD6fh5MK71
iE+arXIM/AbaPHx/304I6aA4zlDy1vL+mq+4yAaaT9G5zKcRiBZagbC5zGij0AWc
LTlbQV7RGVj2uaxETGL8zFRyyzwHWhHEHZvVWcsh4RxmVyfmNsSSIWWIF0ZFMOVT
aZ6PLIxJbzpdLjeGNLXMI004uugef7ItVn9IMod4ve2FLc2tShqyp8OV8pgWCVEh
PooalHwY1VnkNEceSxjHsLzW9soycXz4YoO6cM71TfjWFWGixUj7naB1X8/qeZpK
dWO13SXozCsP0RO/yXb5VqDQk9WjNCZmY1SBtzG2CWRvIPw09Yvsx5Rrt/U6IqOu
2nUGEhibGwTqRxPLU2K1aTKWePzQ7NHTraSgU97UwZOtuucab4W4UnTe30aOKiQv
cwwNzLaC4X5b4wmvLeApQqOQRWBuExhoOAjZE5RFI0QH/1pcBFwzMv4AW+gAEP7p
64miXHtBxVqaKm1tovlbOzzy0VBgoM4ElCI85WDBdjqzZsL+k+WRDg9mTCxqJEs3
vhXE12Z/ec4QQZ46G4lQ1vTGE7lhPrJPtqY2w/DAH70M6vZG8hCLgiGQaCOLH/rE
BxEiILWCQwXdtMDz4y5VqYAjN8l+jDi8l3CxsBrVOYiZ5GAR0jHPTMHq/bUlx1ip
Gf+GrC1je+Exs7BSLxpupAMp8fZMroJACx0UxAaPvEsePtqf1xHLhgCSwD55CjzZ
7dZ/8R6eJ6ZgGsT94osc1xhZ3KL6lUPv1/cZ9KiV3eUVp/RAtuOlTidX96sC3IZd
3ycE6iVF49AzpxULN1wgTdW8QjB7q/CDb0zkfpFFtbRQtVZa1RKD+iwXtQxmMxwe
lCd4lMJ/5TwhEbJZRo7N1hO9ANct8H3QTJcFuF4lSmAw8htdnKwk+jTvptV/DuG3
SMR76jS8KvW6MlqTYCysHFF5EhiC0Ojvd6Zgp9fO41AY1LhdrAR0QryCZ0f6oYMm
I5TLb4qh4B2IG4UNuSDz+jt9cX3S7injUAl1D3tDQBr8ZUs6f4JI2WiLSXaHNECJ
8WrdwhMVDDG+d5wqtwQgrmlprJqZFP2Y98kkPg8qqXuo+VaqbPXUvgzYOH+gF5Rh
AUoUHWE1E+bEXBhEAE4pJLgmwwx3nu3OLCUJ3kjp2gINMdPDy5vSBL775G4MGZKo
0QLjRgP8fmxJcJZoXEkJnnTG9Dt6e9k1DQRVDddsxMNlv8+VoyRXCsjHHBlEFXAb
733jRoF9qnPgLWX/5xPbuZZPK4kgpOW2zvTDsKIcTEBtFkHv8aW1i71BQxX/bCwA
E/yE1hFYIZnpr/Q6IvGKOy+2SMGb9USXHqC1hU2pGiOl2wYXIGFvSer4TwSaaEhJ
XEYAK63ltZeKtUwbeSHkxI2BbmBJRDsKwcrPwrHy0SOsSRvnq3eb82mUfdTGlON0
de04E3iJ1eCrxLE6Dx0HpBVxnOozkC3Y/Zq8TDFs4+aDX3Hp3FnyvFfSYqgc4kVc
U1jskipuTe7poUM7NiS2obrEv46MC+QsjKIr0sdqvpNph1oL+7JfkGg4XwWBbux4
HxjyWAt1K9xyFmRdZlFgClmc7emeZdbcN4FGftedCMxJWqqx8D4kMFX03ttyKHd9
TVSfaFF78pJu2Tt2bv1ZZgsKL99G56eMeVFtUbCv/+vcTucgcCL1tzW+CxxVOw6r
NltC1e0NiwMk4TY5Nqc0x4zdAaVFbk0WFO7EbLR7q5NbhsqgOZcKXcxzrXRFDkrr
TuXV8Px+MSmTMLYFwPZJincnwnc/w3fgeAAefIb5jI/cPBB/bavvcYVC0rnB+2do
ep30qOmVRu+awMPjW5Mbnpv2BzRtk2+S6iVPcWyU8HJGYEUPviwp+OwqFdhSqHRv
Fo8RiItM1/uw/3kN4JAj1p51fsIjcvse6Wo5XYY0Ace71uQktvEix6WzzNAxp7F4
6c5bRbim0rqj8prMp7cewLtH4UYP4MH1NJKWR6fVKPwiNH+qndrys0mhP0urY1t2
efg5egZuOxUF3d04yooeNSdnKiGEN0BY6/CTRxrDFqLyhgngai3r+C4Mb/3i6lZC
GTmCda921ZCrm5l7SaJrbuoM1RK7D2y9i7lJjnIoq8ZOFja9fV+nesfdEx0tGjcq
4yv6VvRjxaOmBcB1wjeG+okVqLWME0k4Rh6msTM1c449DH2NaSdYlD5jg/s69Bxl
7cLWU74UwFYSwKk4eCAU/bmZzvNdAqJwybLOE+nsvuENQpNg6+M1T7TKwurb9bFr
mkb7CF3m+Xhm65lI/aFYWsjjLXvVGliMSEZ8LbGiZ6YUzlGFwsIlucfvVl67w1Nn
KlfjDdQqu/y21rvDWEtNR+hcnRiq0vaQCTbgitjMDVt3y3ZsWjv35HdD1TTYbqp/
vQEt8gxLZMOMz2nc7o8Oq04y794kShBHU6uDCuhUvnhgOFsnNUvMAgUf/fjmpn1O
yh5KX9//7CM/sFoB2MjlbIBFIx4Wa8g15yV7+MxXAjTWf+AHT4Ed1nlebCTYcgsy
m9xZfA9WoaXbjCVAkw91bU8BOreglfhfV0z3+2POhaXHOA5aUDmrSf8qzdTKO2G6
1Fsyrq5GJ7AoHX9cQDHdNEzIVofpP/AH39I66+YQCUKcIgeVopbViZmP75tgWZcI
zWlkmdgq+lXQGCm8DgLqar3GaVrqcW2FDikByL7ypItIwFArja9fEuSkAj7/m1S5
GhAiirtrYSwksU3+OTbXuONT5be/CQPSM4X0IgPsoaDKX7LrnCqITddYINtDqtN8
I6Vq/Dp6W6NyMjFSb/VF1sGTNCUeRUq3Y02f4Fl8XQQRF3fnmrdo3yxdYGsoSOu0
4YXg1RPT89LJt+iQg7MbDQ7dKVGOuTAgxx9WCnEBn/wfthQ/N8gm0p26cVBHkMAP
+fFWCCSi8Vdj8vake9vCNkUiiIxg3cKBfcTIxQn7JzPU21qlWJUXoE2BXn9EnTS2
N5g/TofHskebCwPrUoDMIjCcIIyDxfj9ZlnXVd6qmnPs5jyB6qvo4dp862XlZ2rl
jgA1PyE+lzcN2A3vBaND5RowoxC7qmzwru2/r3ktqT5rG10a2c7GdcjIPvmL3biC
lRToC25xY3tU2ysKxPUj89r5sMyII7SQmM4d068VrBBA7T5ZnAmIKO6rvYF6DCTV
WSxWTPbKUMXQ1UQgUD6iRCP7Cd5JEXaBCSeI+MunR/8IfvbhMcJBXCgGuRfQzusy
mfwBLF4RQxAtN0l0mzG+BdINHSVyYB9hIHiDZkXEEkgmjtuAD/Qqr5J6HcmTcSGf
Jt2EnfC6Vxg/gn+j/2mZOitO+mrKV1g49hFb2pJRO4swZQ9YBtkqn0NxYdw7kk51
Sjo0lAE+DUb2f8hhRz2/eBXNGUcNBIu95IZcBuhPLYWypBLv1xfU5vOVd+618tFl
Ipl4FjKUM5Cehs9PtYPdm05IoXCAM+smAR/jLiQNn9aLKD6O3+bvOW4AVgt952Ho
0BN/WeHYOTVIPfcJoDoJ9lheJde7NBxa3zhiI9o30tDOjvkSTAqwjMnwKObuxo/D
cfyd8t9XeHCoKHAT2gLaFQQlcLXlCF6bDK+38rIPJqoVBUV2IqGHktCViumBEY1L
+unC10Z5rbwUJ3Rzw5Odmco+gpOvlgCvtF0v0Fd93NvW7w+UkS2Zf7X6XOu7Qgnr
1n1UsFlj41uc8kpdhN9b9McL6uYkpOE/yy90oUfBgaWQ41+EWGuwinYXvSVAsJEj
QwDSSYsEsS0RhhhPqvXR1Kcah2SKWox9rzyfeVThrcUuJjuk5vMnnUt/lN7MS+p/
dbm+L8vhJh+0LNMGgQMwPZKyc5HfFPYf/aBDFr3s2m1jGCzD4JWt3UTBDnSiufEq
prOR2YF7yCzWfdswEsBNiECV4Dc6v76llRT56sBz+c4gG6JHfA+DbC5nvMb2Hyd5
wDGFvFZwYj+Sn96MEFzE9WKF7OUFsyv3qQtsNooVLPjuh9cWElmtlYE3NT6DhuVi
qJtMQ8PuArQBedC8NOJ/9rxDFHYF37out8epvSYmCgFAa5Bd16KCtycUwHv5jZPj
R2bQjsrLnodHu7kpAPguRsDwS0KNEDJVdH7qEK+UE84t6hEbZgBtidxdIqAP0M12
besWp4Oi2sM57hcIeIxEAbinxY0QEE24iws6Ha1Sq0xnTYp1GrhKYV+E/YvLAf1A
QUG1OSccHnnthSDMFo3U4Bgds6DERzE/WjTahJbbJ5NjBgeE1XBaJV4DnfMG+UPQ
FCQltqFcqlZUWR7JaFMi+5xGN7cqKkGTkjZ8nUbpaPQn44G+elU/Zay0vyX1/22j
qqk9XnXPY1enl5Eb0UWw82U889foPbwMxFBIJb5MrOU+5d8p4S/ec+0ZnqKiOIjK
jpe4bdmoggXuKVJjGOlFTC/CbRgkM+b/HE92kTbq7DmqLirEHI9cCEWstKeOEYlu
x5/gVUMD4XD7nhp6atAqL2O4M+T0X2icAkY4wKijtt6jl4slLzjcgx9eRLOmmsjh
vbxrt6mpSs5SQ6/cNf8zHflCL8A8WpfQ+ohsjHv2VkkUPv7havnLk6b+e3tUVm/8
tCLRCeFWdoALyftgdV4ucyjkMz7hUEeTIyyYHYnmsdnxlAR6k/UkjhRaod6ybnqG
4G2lXMMFrfX88VKE19qnBWV+k4P4T6fTfd/Yew+WkUTIcKNVi9XllQ/B25jKCWD0
n0mQiPfuU6al2nC/1acneRn30TgeP/ab3sIRoDGJCukxpnUzXBq1/6YJupZRFLz5
z61Nr4cxiHQabFruL7UxYnWEOs3uhobSJkNKoNh34ns7SRGbQ/vdj0bSe0dkZyJo
sIXM/7yrDTO0FzHbmVRC4I2i0NPjuleKJB/6b6NW/KtCgdnlRX1bGxO9mP+lEGWq
dtvpjEzCSRaPp75ib2tUDLIqhSJYgFxsVG3aM7tVBkPJhIKKY49o1AF+Ur57ubTm
LCqAJSuH68XGESK048YvuV/1W43T1Xu5GgVWYMb4nj5IgxCDItFNHvKGR+ev05rO
w77Ey/6RXG8oY7zKrxcIHThZvm+gDuTJRSwdUnpY5LwnLnteEbU7lTzgcq6hN3y3
vcovUllTu7SChX6e8YN2jxNd8wV3D9Hbw59PIUh20bYOkFVYpYuvF+qr9Xbbnh0Y
Ps3mQGYTi3QSLqikJV5UuO09fUF8/qFDuBzilt3YJ+bQMFYZ0bodKo5EOPubjJpa
0FeWwuMbqiUokImAXdXDREKQ/eJgm3sXVRCzZEZQYMHejZ66Xb+MRusvOlKai9Dj
BCJVJS4oR8cphCxaWncn1OBlt7YhNpW7FidpIkS38K5wegCK+fIaZE6RiHHkdZLE
LCRSaMx18wKDvNa/bgnxbSuEroUN8cOClhTPQl+qpA4w4nuxAY4SbOFlv/nb8KkI
eLyP+lmQcs6c2RGsvdNy7hSDBj5XRAuuKLEwqUHa482Mrxa8R0nSWvQQ4Byx8NRy
WtxUWT6jWXNdQ+TAh82OM7xuMa8teTUz4fmjXhinF8yq7IcHa4/EQAzYIrDqbFfi
b74OJskiH34v4o8dFod477BYoClrBbyBMJ/tDMGBKE5gbnvvfFM03W4mgLDAnKBr
2dlge+egoh59rzAtwWo3fnmG+k/ojQMTKKCxyoSJj6/DonDW4JzHvfH9S0ZgoHFs
vqIlOKd95cqDIZLhclaU+ULuOtxlefZom+vxxnlEyzOGuKtqOsTaVJdilJtvEsMx
4MXhm1kbo9gdQGCFY64VM47vnQ9QAETa2eheFKCjccg5IbgYgsU/XddsPEX3A3SJ
AOGXMm/Qis8rtuEt0uE+WYGwGUVIkPvlCpHIMu4H0OHyzjETJAJgGRhd0Esdrhdx
Pod5TWhhnnblijDcgb6NI54M7wkr6UNzqcQ7mtacfRPYJkfbVrm0gejkA1qUUFk8
K5jaElU/5+vdzTubkW8DnbXKB4W1Z6hp3lRfWa/SR1EDL4BNZFMN4+ZNYN8HyDd2
LfA61RcHZz5Xlhem2yD2j+cx4Xb8rZnBbvlcf9sWUG7pghCm3mnHLw7ahBhnU16o
3R2TuZdEdRmvkP5WeF6oVvX+wPaVBeanImw4cEBakw4UB8ruTGmP1Rwee5AdMLDL
kRJJXl4xMv2uclhrG6AawrLUce43Me7bZiuHgLCC+62WV9n5jLOkXXsKj+zR95LW
DvjmwrgHW6z8IjgAFxEDughI2cwH2rS5j5cT0eAx5pXPZcYR3gIIO4Ev35zPHsN/
xr+LOzI9EQhbFBnnAv8g7j+bkMmjkkonH5m1EJ00ikT6GmgX6sY9BZjDGKGNpHyn
H0YLQemZZzwWsDijG2RyGg7wC1BVFFNIhP7kTCG+i+RAUCn/qYBTDNV60aFkHeD0
f1biA9h6HHRhA2aEWlOcc5LP+N6EMB5s6o5oFKl8xVZ4r5PVcMdxUSHAmi4Mw+Av
b+my21WFwWFt4EWoKyFpp+9clmGbvc6A1MWfHq5brRpAgoRstut6UW94q7S6gnW2
bwpsGoTuwZAa6PVpi58xfXAWdARtr3kkX7G7VDURCKdLZOpAhKef/RV8ZM9c4G+F
jk6CkYOP6TeETEgF9VoAnWfhjjDSbpPqyd/vHGciD5dtkpeUYt1YPTo+Yu5nGE6V
JXN1FqKWHWwctDYe9rx63LAnVGgcBT+S4u5lbSHIpudS8mLeqphXCIfTTgeSlyEn
sJ1elsUtDRRn5OdugATMT7pxMd+mUJ4EQj4lvBSORjZTIyYnX7YssH8TYc7ySaNC
ybIdhtEStAFf9FVju8iMCK7TzmKIiGhvG5Jf1Gf982fSaOGOoXPoxT7VBMlkhsRv
lOkKDDfjns9FrsJvszes6HnEJS7vzf+7mL7Eo3sdGwGJi09vntixj+nV/YFRvYlt
qGxCsHyHu0cdkEa+FDwk6W5SgFQUtfUKXMe1qNYEnpzLKIetrLZde7Ag4wC9pswW
84sS3+/q8SL6oBZGn3eXKEMyUl5Gc7LcwsjE8lE4zYfDow5mPMcytLM8nQygsDXX
mes3ubyisyqimxm9/Vuq2mj1F2SVCDON97z1pA8+5cVjLqlnNxueAx2XaCs0nkJC
kSb1sb83skYvywdWmo0/V3lZ/sPLvD3qKVLIhWZEuc1+BsM5+Pvw2DgH2iOEdWFA
K9w9y8ARDM5KX/qwlNVaJcGMai29tMjy1Uzv9IGPlxRMyZhPcLlOEOdr9QvoOhwg
6eswEgaVct+ZJ/u2Wgtma/fsvAqnO6gAWPlG9WRJ5LYAdlPhfXlFabbtPEc7QZe9
xqXrvys44Ex2RBFOb6wV6gsCdPXFIHdOsBQhD4O376XkmnkRUqVQc3JgZ/AMXBgs
lHuPEjQtQ7g82TG+0FyyHdqYUNhTKSTd4BqzcblO/JHtM74jr9U8WWggWEdSvOQD
wRjFVcdyUzYdz8rPdzlQiTl9l9MPocFraH5RCh7FJktqq28zmo39jmme8VF/2fFU
iYGcTRWTOzkoxF9pYKqT2v/3E2a72OyRQveSI2egN6FpuaqkzuZRtTyfqEIIt8eh
216sR7EakHS6x+qriyzuVRCBkpdQUhWTRnp3FXan1SUkReA+oIR6IRlv33ve7W/i
E1SnVBK9k4sp9nPu8BGYXaTgNfTHNOM2oodizZQmne28FVQ4qzk4TsPY2wdVQku1
+Ub7YAgEi7UXD3EMK3rt2iYs1G//NwnucNTZ6QsUPrD+xtiWi8hfeU5uZuGF13yG
vCxeKxoHtuhIjB9ryUwQ6k0LNHlfb9f7B81DVf8USbrAtLrsb5yFIEZK8EY9fue1
rrp9K3Eh9MjFB7Sre7xrrk+G3xRpYPbaaBSuUhjrND+Cc05Vu1g+n+V92v+D7s2d
ypZggFjfJnhgK/SdIwfSDPTyFaL2ibcIzalQM52RQf3egbbCeJLtdvjKAcgBg1jm
ZILhCu9S4EfPqU1BSzSlu9QePyd1h9koJBEvMdqBJeos/JItXpA5iFO3cV3s3I3F
4KZaCJU5UaUq3Wq00RZ8Ei2NrK1r9Zwa+Ok5zlzv/COGO8LMjN8FUWWMGvbty4Fl
nrVGVP2ZxVmDyqHbFCI1M9CsZ0IT/JZkPzGP30xyziJ/1xQvjgg/rW2YEv/q2HTp
8YjyhFVkeJsfgZly3exvcC4kgOr6+LiRJZj2XMxgqEFDHZzFun7h0JaLTPyzaedq
4TFDy1Da4gJuZkCJzY6ZYI0AdxK6AjoolF+r4axzM4MQCdTI5k6lu0rU1nX5qaTc
Jjp+hr1pmFAuXTqVi/k6TCepYSMnN1x5FWGNyeEYBqYayehdkomlneUqr07eVRyt
Mt4Z7wjjmPdSUXrdBQ0TUyFV2ZFvwfNmZeTWVX8X1sBGFcO9rdAzHXddBXtv9GP6
HB6oeu33Ek1+kcQzyqIlX2V6hspKTxlCHS+qPmDj+dIDpqpkQt/35y7oGkP0CB8g
MQRtId1UI4pCAlpmQNtFtV3sdNzddxqeZpubNkF3kcZFgWkHT/YyjfxWpzmQ4P3I
AAQJhfXUNN4ZJJ5c7d9hbhmpSU8UJ0URLrixu3A6ZBPsqVyC09gG54vdYS1BobUU
YqRZJCvxqgla3GSBPQ2ukk6SMKZtl9zlB5yJkVtODkBgufZKm0mXDt6qGq5RzwjR
41YWgJH9GGGW+czkEbAIup+KSbyc6qXvfBMJp/jsEfcZjyOvaRW8LdQ6PC3+vZCa
kzkQYdH/Wot5G2YM7P+nc1Y6Jg4a5HifWq2532jnQupWgsHNl+lXJ2nnVUqCOhgF
rElVDe0gRSKbUE6xgDH5ER7FuuKG7Fdc+E23X/qMkj/BSYX1EtiV+8uHXMm7cHFb
bpuNYuSSGeDtZmbYhsIdHUIRt1V7Fgjfc5KfEorcCUTJ4aJPGMvOYc/GoG7ju9Gk
nngvjT9LAeQRHpnt8NWI2pOyePi8xkZDZSTmF8xY1Hk5AY1jKOxTzBzELExCVtJC
zgQDmLtrLKkv3xvfO2qPgSdiJdSdSMHelsm2r0R8YiJqlyptKlR0f3g7hYfO7DEH
4SnrSIrIkiRtLuwdJyPU4Qjgp+N3lO46V4Y72Gpk0pjA8qUyMURXW898nAR40j4z
xyvFb/VwDak//zzRI4jquDnHcPp0p/FPznjlv3tO7+HjvbIO3McrGY/ztSUSmreW
Bd4Jy1PuNMTIZWLDSXPIUYetMTQ+CbMEce7x56fZewVjeZzgOXwo7n2VY3Vt5gGx
n7Gy6zn8gR2Rr8EI9SeUjL/LCekIcK4es8JldJBmfTIa4LQU+j75S/XxdNEb3pJd
vBvmE1JzYWdoTMslHxKa6h7ZAxvyq1Ndih5InEbWZxaMcgf1iFq4MjuNqaz2kWXC
eBZlKhTsF5z0WbtUT9WtR/PMpO11lQvs4IRJFwLvn/zaTJ0eQOG+m7Y/1U1zchdE
ItI84vjT7iTJXhM+K+/Oi+pKpNaQeEx0eKqK22+oh2T/gHHUnP5mzjcbp9pAb/yC
sxbyN+sWc9tQE+Xs1/1P2tf1xEFsi/Q/82+NTnWWAAvuDAfH26366HeMqO94/XXP
va2/VNwKO2s9UjbPZz67mcLMsEbQ/e7zX1hwvEXX6ZAS+y3scW0ecJygQOwoCMnF
9TCjsjMHCqJJjZMvrfWrWp5LpjPHBxVYtYCrLWTnZn0AT0jh6ZFcYiDpnDkKCYS+
kxhDovss6IKUDXp4AlKy9z57cwlFpjStYZx6GvKHLOzSOqLwyet9To5NEknYhYE7
+4H7YZQ0VXchxCsG3RIK0Py25nuBldXCIJucN3r/qg3pIFqGR+G5GyoM0VLCLpy0
rM5GMS7/9ht+d4e/hid4VJNQaF9QB7yp5C8Q7yLtDaJqYdQS4AOKORp/bMWBOOzm
qoyq0vnG5ozVXL5AYS3QtY2UuzOZpwVZFz17QXpAsh0VeVgdIAI7fkbO1hNFELI8
Cagc7fdhiHCohltJXyse5tygiggkQ/zT/2Bvsew4GwPDqZEzrrwp9zICfY4WRqTs
3wS4HPMcJaofgt7Wv1cfBuAQks12gJft3ArW7v2gwc8X6RdgGzWQiIVy44VtEr1p
jCtFtXyKJQC5/gFsznXcocR299uXqwf2eLf75YME36uYv9u6w/2E63AqMumM0uEG
kNHS0DPUVOnezfDrZ22xAue3dseLDdiLXScakzqhSynPWDlvLnVHzvjMuiJC0GDn
l4I2trun85ObycS78gfzUalvnc0rmPIWZUGOHSoP5k6YHM/9B2NdirTf+fqtsyRl
1yKKV1kwZvuMWUkQvttwABFlBVY2A5YqAqZ613C+ngtkTWUjoRxxQ7nrJCPhrVR3
PdnPvh/uYAaj+75RPC2gw328vHHMv4Eg7UXgZJv5OON1SgpmLPCJR46Z+r9kp1YM
6gjMHiHmhj8F2bCtusnpt/y1caUcc6J2Zjd+O6dcNgOuGNS3qQcAwNxWQZ2Quu3r
DgmsAMN1gZZkXhB6yyt3G3XvajNFuwAcB0GDWgU1Giqp87GzKVMnKG23qMh7R40F
l0E+1tE5kzn/JWcEjq61+yb3N0Qs3kTQi0ZlQfRozsWWqtar9aVwojYaGNRHhpeO
0dm9AIN7iRL5vrqzL1yLhV3AWuRgAM3igHNP1gN6NBuY2aBNopXYyE9wfictWaoJ
gJoB5WXWGkX+c1GkvY/wtu3r/9GrJ/FNDRu5n1WtEQNFaHai32AoIiQaOCQpJLZN
pFs7En9UZDv/XUTwzV2mPR6DZ6IaJGdJJiGCHMrebjNPujuHShXpHNCJ421Ga6EJ
oN86rolz7SG3WZTnGMXoNkpI3sNAh/YSyRdXnU0lnPkXwSC18w1ROMebZzxnzfNU
LjBHJSqME9EmGR9jOIgsCZN2waXBpRiBYaHvinlc+x6zyfp/UZaZ/Tj2JtBohIpw
dhbuctCCAyjFSE4EFzuB+Ohmy1dgtBNogLMIBr8Exq2aeZsR6tP4q7F0CAHeaKlT
AvgsNbq2lt9YpUOcjJv817o5DNgj17+Qj1tvkwlP6qt6i64Y8YgZBJa/ut0rA9Vq
6sZazpOSt0TWEg138sJd+rnAoElPKKH5F5HJakn0fyIdX9ed5Cnat7DJOgG1jExv
1gIB1ukQy1Rg36LhPJp5MFAHb0e98v3efvbGjSq+sFWOj46IXwANrv9ZT5ibXS95
QJjeuGvoyBlm+QtkkzKAibZ8Id+MjkgfOPh3dI3lKyzpsRyWycStZRJIjlBjcARj
lRBEQB0ICQ8mp1EAaVkViE2sgdreBlVgqkzyFZ/6Wgm7hXOxJfM/KYTcFgZVYc5N
j5BA/5FOI0XDD6jBsDi0wsg2UhBeup0m8EpC9+6OSlapD4GmkNRF654L8iXHktRT
We55jqHfQI2QVNufXmwS4706Fa3k7K71O+sfhWq/fdBIGmWS9J+l/MasTN5dBaaN
55HkJTWV9L5U5cKgKU6gMuxmu8h8Bs1LZBgDOTKXf4Lm5pMjaR5tYiwIzDy6XgWf
kV9j/6Kg+prIAXfFmvm5e819/BS58UCs4JUbA0Ef65ujoSGB7CWQv63S6Rq9Px2X
YjRMO2u66QizVwdUu5yYwQsLdNigASBXrmm3/dMpDdhlWt0dtjB3WCs87uALpgb3
hPvkAFWqiI/YQxKVQ0MFHnm+Acfb9JUQ1I/7YUCQv4R86SJGYPzUncy4xnCL/ff5
3uFtSINh06kTmUuVCEYE69w9wsztaoMbWb3fXhNej8coORGCxfGhHSsE1nq7LCvK
WcuGsjP0V0nEHRN32Fsx6cKwptfhCb2ibLFMJfFCnqZnHEpckcxYG5hAJvHArG9N
uFP1SLLJhdPV6UcxIEogL6n9hpRgVc521KLGWrkcIVg6CYfJqWe2iFt1ulGfowLF
x5j0yRvWIarTduifMwtZ2U8DmvtChHZnIog0jjXxfKNTPY0CIAqrfcem8/IS2h2/
/6Z48hOrDQ4oB8zdirqOQfrclnT0qAzcCXzhIlD2bWiR7a3lmn2+Z7cVF+as/NST
mP5a9P65/vL1eFJkE/qTqAmhadt/alIdOWApdFifL1TERMUAAjz5TUWJozr2TT/o
2x64Fs1uk2snL8Jr45CwHCGSICyceWgJ72N+8xZDO/I7gxDunpspNaorBwPAZWgH
1ftR4kLtt1rhA8jkY14dvo6h2M1wqE2Zz5mZFuhrFlkWU/qsuCUib3F0tj2GvDP/
EE2amtFCT5nxXF5VW9hF+4MH5tTOZZNg77p+PPeZSnlskgOH2hVf0Z3WnOvvzMzc
hRYagLrr3G8I/sW8vbus06vE6fCyMYUjYw51hpvC8qvvkU3uYNdI590sZ1VEfoRT
ZudIhaNAek1TbTgcsqgFdSgPa74Dvqjyw1KIatvD3nS3h8nMPt0y9ajl7B91jUoV
Gh46pnIWVwlwEkyV9YIE+5sr6nCFKX80ZBPl4L+orbKV91rQR8aswuRSJTtMfKgl
51+n8HVet1eOgtIg9QNrFdng9KW5lF6B9PAq26o1DXvg1vhFSGRPIAkfdFAuRrl5
QjDfCvPzJ9lWiSufLwE+DwA/BLw2ro/Et70fj706EZx62dqAXP4bGgb9av7fEsxs
J9qtjbLhQf91meIQbKPc5iN8JyF1DSfWDhkSDwdKM5iMT3roCC6+gk/B0zKa82Kh
Yhu9qNmz7tuagxa5DizsFzZbG1i+GieBLHIDk9n1pZde2VCFLt0wHBA4PbyFjQCh
xIslKtKWtBotN/eYPWFPYdsLm4cOQwTYi7U9ZqzmRBzB5jPjk1geXtAMSqamQKk2
Y3E0tua9/+cgknHulI7qjh30oorX+I+IYDuixLT12U10rJHFJscsBpINJh+RQO+L
3gjATVDf6t/KG03hCk1pAtopHWQ6AZ+6VDHUoqKSAsICnZCmC2v25zzBSjGky0h9
jIJhJmQrvhrtwYjZmVzSSP7Y6/tcnrxFj6iZMaB7f+3SFxApw1pFdOhy8N/ZpVOG
hWF2afMGx1NtA93UrvXqKfWvLkplMZ2BrOYOcZGto5F9CJaVyjkO85EyOb4JCJRW
ahuym0FyO4EGI84w7iDyml58cew6fxbBiu7s5Z+zFcqT2zlRZWaAXyH+PRRJuHcb
XXakekv8VEN6f4fszJIBxT+PMvHFxTdRSQSCfoAaSrFzfggd9Tp7mBg33PitEgzS
ksXI1TV/tf1Kj8kkasM3M3OL4olDRGfJTfcuH9vgEdGya3FX2/0zVAG8+oTK4my1
6kn1xhn9xpLdlhwcg8TcrNd+SJAjP2toNxRFivKnjtU538RMjLwSQMsi0Ss68OPT
Sw5cw/Ng5NAa/XQelDP4M9AyHc11KQBpDoFjDoEUkFGJu73s1/QMUcs41bvsjQv3
0/Ly1EKWTrW62TkvIc9tc/IYBcVBPtGDoRz2eiRIHI4aL2Gtc4hTaPa9IEDg7Tum
xnbI4hlDWC1j+nqgaGaIwP6BpsPbNsCT8CElvRX2/BfHJ4YAdhJaJJGyOOCutjhy
3nPTW5tG688nok0GydcgOBcTuLq1qW3jS0iRYDBmRnpmZmu66Q2d1BEhahTlsebN
/O3eiuNuLl4A39jvwqJ+Gmja5430TvkYMeS+s4lvFqn+KyPC+Od5FF5Oc6LY1MKn
6R/0M8DR5zhBd8DcOVzJWXmtt6fJWQmbByts8F0TpJCgE8oI7nfAmp/8RNASDBk+
8BmBXse/5GinZldbUZROw9WnDzd7aJwZ5WUInxrYehTDjpK3FJKZmvZVB6GHZJD6
c7KW1X0uToS1CAP1+knjC+n3e8XU4Ehpo/yS5DtR/mcWVCUQgBN7BrZdAi4BmcUw
/WqORwJu/VSMMfArqB+z3gbbc4ljD5dFKoIwjPS3+472yVhBiIQN0CnkiHwhS4Fn
flw6KOSf1OdngQP/9ZqgBwud3n3AXBOSb2DmDsQI820HILg6A2EfZr0wChbIaFf0
xGcAdPTNCAVdYnSrOJmt1xHx57V5bObxvE/MrGos9DAYefejDNsVJh7U4ZuYOIbI
I59jU57Fxsb/YvZ6RwTaeqK39zHLPj1Tg1TFYvtR+KpJv3v0TNc593DCoOMRsWSh
RzQnRa7Gi/Y/33VOljSZARjo4Njf8hzrpz9RhQIRoxVpauLU9Mwea5xuH6jPwnoD
IRelaHtMNUUSuUwTc28B5tT3v8usdxiOK/ptVOn9EN4R6+G2M/NsbSvMX6M3mGbb
C8YK8poWzao9s7z2K9lRXlLPGBGck4Glrj2dD7VgRdfz8gJ4ljJXdQMk//gNsGV8
pdLFOYExSeaaV10l6f+HEAY3Dj5ZCNP6NrWXq9B/QNxLbcYVor3b/zwsoxJ6tAfg
7fQfx1z10C66t+7o6eALvc7vScqWYV+MCVXJFnvEhNCCDOKBzbbWIokQN2MyiHYr
NAOy0z09XUEhteVaqmSdNQMnEsLd88cCfsI23Nf6XYyCinBqIl2bxRY9FvIRWCdw
Y7ESdcKyhYA+fhkqSuUUpWI4MZAYTvD9J/hlCSnRrRN+O7R9TCDollGhLgyalDv6
DEoTXaX//+7HOYx45K3gOD3myyRkuMvZN3niXMbkYvnXQrcDX03RV0tUESzRaIMh
bwAQ4BEVse7ta7VHMHxHmrCi/rMihYyhzA/l7rBGH1WIMQCADPVqF6SDTNPHA1r7
yIC5NzwEdKS60ZYn2syHIrZSJS939udU0vHkHkBBhAkW088icb+1bWRgwTOaO7OI
db7it9ZEixokqS4RRh2Gb5zRmknubG5Wvl9Vqow3tEK3BoG6BBgtNP+TkfPgbWvL
R1sHEnx7IXMyW9vFmvdvpgj3lpBCIxH4dNvzfOun6FwqKgFQ4QB0UyfaiaILrXMr
vBuVz/Y5cMeKwVzLpIz85PDCzhVU/BghN7/nT+EjL+BtIaMaoZx2tm3LLbmUPXa8
iYxim+GUCJ/sma3ytDFUhBs7wj03raU4dTEOMTYayZgzrtPsRPu97QjZkcS9f9j1
/Jc5IB73gANG8VXTE5YJD7VjIASN/F0TOIG/7nmQfYWd1P73XG6ImMR6c2t/+5cm
ZfPjbpHBOAt5wgpVpHLQhshflr2Q4TiI4AwRZl/3hOnYD63jQi9bMiJq7r4044GY
PUgb5Eba0NcOO1pJj8nl+9fzp4H4mEssH1e0a26Ki+02OL1W2RmqAPQR9cmZxaSu
zWIUfv0t/J5zQhj4wtId3RznuaGjnHgNgzwMsRzILgu6wNNCD6fkI+GHNeNt418j
tYexffdPj2bjquhvOkK9couit93gGhF4Nm4bgkehP+ZhtVuTT8TWvwOYMAiH3YTK
VnRFl6vla8WHEEebNLLT6hmxck5hrJLnnCfhF58l3Rg2b3aQnak5pvIbbjUSzPep
g/E0tnnNmimUUpUSZToRyR7ihoXgYNwrFqMU4EPY7BVkn8C0nhcQTR3tqUN0EnH3
WutaIGHw1ODMHmgLr83X7NWS4dkJMFbV4uZnTgb5bYGTc0FNftEGVXImud1R6vDZ
fKve306C0ybrB2UBIIEmUy2E75a+7usXpCc+iGFgtGPp6XcyPtGg2GN5/ZrVmLkE
Z+I1qLrbTtDObt0rIu4gr3Y2xHLWU527V1kTeGwfKFbiw1NYIxilmm9JjQh/GD+y
mRNUKgbXp0q6gqFb5Cyti+3ZTGd0BtQnhm7wMp1PQ59aEtxGdOCK/COTY691kybU
IzA2SCh7aL6y9Dq7WS1qZs1KIN4Ojwn+dU8eIQnJwDT6r3uEHtNoe6Ts+l08t9x2
C/LwuLxbG2Zv8k413dFlbZtm2nAMMFDP6R4RfWZE0czmhrPRqSac75PCD7v10q/j
8twVFWoBF5dT6qPheV2sQ8rOz1smdr6IKTg/hU4TCPRH3+5hMQbmiB+lrigjYV9Z
KFQ2mrw7OAPjtGVnj2maaiwijUKyJTLtWVilWpD3KAFuyAqO0kXxLZcKhOt1ATSq
R1qydLCbauipRCIbUQo18Z06NLmJfJ5mBzSA96mGZTLi8/nxGMQMolDDj9rRuBFs
yA6oAuyvMOl/1yse/998LZ484ab46duAlicpAuWohxnm5eOm2GnblrevRBg44Kse
MaYsbCGYkyQmZ57LKHdrCvv+9q5JKJt4x3ZIc2Ehj5Bbu2co4JTTEXZ5OwKDQbJX
bj1oWSk7W7QmJCSDiixQFhggcUPOW4xOA/mbyBm92LQSnYpUPi7DFGIRSIO//U/T
mHvzA9sCUuAiboB+y5JeC0UWV8I/ap3MHc3ajjNf6AQqbY8qwddYbF7wdyYEYJJ2
T3SmEbMG1lXjnw5M8jdSOi+HGPgp9BUXEXnWMsEngrfiOtpiqf+lJjkF3xJe6HrL
8r3Bb868WrS2KZJXprQ/Ue7yjJoOHSLmZH//aRMFUU8eQRxRhaafyCsmjE0imZx7
mINqsfCXRP4J+R3D/tNi2uLLMy63ipBpKyozCO5VuovkuQFH9SvXYdwapWuhtj5N
3uAPdC4WgAP2twZ+Y7AtOxybBvAYjgsqD/Q+FFeBVuKOzBYD9eYKi974EaAK0BTN
7VfSodF/MhnUTYSFp6C4At16CeWVY7EQTSSX4t8mO9MKMv85bdcYamu/eDkw9otc
omrLiawCzKq0wOh0OOWQGcM5meMqPxp4PzPxJlSk4NEUBR8IymHHf+k1P7x2KiP2
/13dUvbr1D6paLHxi0e3qQtMm217C/+PM5Pj5SORIFRS/oXYTfiONI74rq/KeeKv
5FBvUfsXzoLi4uKIT8mcXqPZNHL5HJ44wtLH8fcn8PfbAVP/OytVmZxRf6Z1zMLi
dzu/mhdkO+XXpjznpz0sQs0tMPKExdpkHURAHIjAii/0iOZPYQU0N4BaVxVc6+im
z/7B9SD+fdn4kx08UVsfsrBQGTgKZGIzslOIf0AMPjA/T2XanDtDapOKWO40/8wN
xQNmZqStnS16LRpUNtTqQwuspIbWLsWK3iJqggF+8KXmQQQmq9GffqhVNDYMx1Ff
I+cgOe7SNWtBZCi8eQ1GDvJh4g18ERH8ktv/KDHb1/Im2O5utIMTWTv3h/6vVUF7
6xyBgcV78MWZbgac+109lqezMiKXfsb+XyCQkPef3/fK0tEfs6Arv433BVqaPiCo
YKDHxDslIfSu2Pba6M8bT2LZoq5Kpe2N0bUhntmyelPh1fNvylXQha0SUHOjJkBP
ufloBm0PcCo49QyQ0FERK9z+A+dIH1KaVBFUzwj6qZxXRlCBz5CU23ZN6iNdbThz
S+5ot/qFAkhwksPyMwnfrM2NyasUwl+l/cwmZNT8ilr1uE7LYr4VZ7RATMmUTw6+
c37C8ob5dpeeMahlpvWkUCFxNdm1WOR3JN5I5XRrE90psw6Ddt53/2lbK/Mawtxm
dLuL1OXFzMP1Su6XzAvNMQki+1UrV/xyrxHD3xxBQTgu7n7Xw7QNUVyr7TxYg3Uf
EIfHcmnht9DoIEj6+rZxolilauznKcuko/5i+yA/pL8L3aMBNxo162lYApRvGqr6
uFwwFaiIAS6kUJx4uHxDx1v/rb7xak3nHnNmzEtBwZtgeQXtgGJOZ8Uj7EfwqoLL
iRnPXzegirpbX4cVy92n0gaftqEdlJuARgjEs7AjPcxSs9kN9wN7599mJRXIo03k
CUsTzrecomy9N/AnMpG4MG2rfJQnvB/7kQp/cj5euWImUwkubLeoAInCjUEbb4zh
QGriJ0X0IpOlwOqBa7PjVPvorOX0U2gS7mn9YDXP/tgXbgLk6AdoJP5OzNK61Tar
5gPwbjLPQ/ejvQvJFX7UTwKjl6qO0xNL/Q/0Oi5BJcB4x/akPMxqq3VAlVMNdoY9
Z5jsRhDBcDuRSYNuV7lQDC1OAICvhuwYf2I+aP0w/p9490j0YFr8xf7QV+9wDmMU
tY7NzY44M6cmioFH5hYAzbIArKBgdicnbmVuzjOiSVbg8T9m9e/vCXW3FvY4Sxr8
orLORmw6BlhJ0cDNi1QyyCVSPxXqMdR1oCU2htQ464ErHQWcwpTLYWbrkE4BdzLE
1cslaHqSzCQjSlt0YHrmL3YanwVy61gM80PmAeAlQMmvB07asgz/AtghxGmyZWDY
lw5PM9P8UDsSa1bZEh27nQXX9bgphZbt4p0Qn5M4AtTv4N/poWFRt+olxxKxXagn
qVABw588QWaHas/y5yow68KqjZykryWOF4A70tzjdB1QPxj7bUEMvQ3T3BxJMzgF
CPViBQ0rtjish8Xsc0Dny0CeuyxfQfIuR/ouYM9BqPzQ84IWiKYtuy7GfX50nH7w
LscjyK2j7cJiY8g0NqoSFLTrWN/9JYAhxJBNaE6gsCk5UC6dK4AWHXxdfdvZtAYY
blYFFcUEdYktSa+ZPA4XrmVZTkYe+cnvmorAM1fQiMMMhnXFATDQFJ+qOHnjQG0g
U4ilyRTTjFC0I/FsiJjWTIPIuZRn09lHzgRmSITVJPrn7d0GONFeodVnct369WMC
JqKy6DkgLObViUgaO05imvVhZV1K2WswLP4tvn7FUMiebaA+yrBRN+JyZ3skHlWW
TDLXk10xJOgn3WvdIE6oCqvkRPutR47u+khBzsCwcqPgUuVplyiFA9F/h1WfyISO
XdLznZhPeU+MmA/yte6BHRfRTjuLI6S7w1a148tCg8QoHzgf2au8K2Ybj7/HayoN
d1t4hp7eSDVInOrn7prwS4nBK5v6FQIgXMLV9Jhpq57+wC6AnDz5V5ieNWapfDP3
IWr7vvpUXGlmguu9eOor6n6u1zR0lcPVngNdxkQq5WdwgpDKlmS2lizrjym5iMDJ
QEms3/KvQsTpoTGy2rrAFecfvJFQ5a5gedY6oR3e4VE5a4e3OehLmLEdKO8ph45B
4nMZ9sVDTnMP4atENR5h34hN+gB8z4LF7k5tHTk/GcLC4WMzbtUQHyRSx5z4DYba
HFr1xcK2Rhh430eHheshze8jef/PR2DNNBjI6fQGDER5hq1HLmEHqlmarJyBc3dW
G20vv8uVQvH6zc7Y6CojBaxqnmlrp0Oa9nFP+YCcGFSBUvuFSEfksiPlqM7muFMK
m4UqNwbQk/P31KAMpZWXFOaqcgK5pQgSvWuW9E9c80iOzcLbeXPaOgqcJ/gX10uV
PX0+NMbTxnzbfwd+IPpfFWG0Jnw44SmC0rs/4q2QzSdqzgjCgP0STLgtNbV+vuI0
KrppsGL+aKPQsOVz+p6pqnGmApHbKV9w5vihRpsMA3+yL59+1aoLV0Yy2w3qD1A0
3JBnMGoJmS0IxRP/+d5KBqYn8CEMtabeqDroRwGfvowMxrziqVIW8vs7L5041TjV
trbgX88ZTjJY9NZL8gzmG8F5RFOHjLwhVVWMC8F7bFK1yZuY3/RROlc/hT9h6JoU
hg8TTgS8tCA+t8jV9jyCx228yuBSi6/UDPMJzdyA0opJP3aQyyWMH7xmUWxZjezr
wKKk3/+HMnLehqt02IQFBO0lpqbKH7/DRlBy01E8XoccLHVPM2oHsR75ftAEAYq0
d4iJPLtJoUlWp9oZv1IwA0qfRgYklAPdS0yFgreTFr+3/BAfkcG9efME/i430hc5
NOhsN0EY9vOPSxf6/l5JDv3l7lEyeuKxpnbMpCmE0RlL3TD2aGjAm5aOTVQvZjV6
8ESTrbjEzy838eCsRx4Hv6j60aGO/2+fY3KDVVX83vLeeIa5D0IQQsdHZT5Osq05
x1sr+Ns/NT7s7hqSDykOIcC2pUvDylJV6I/GotDEQG41ea1Ro+pEbQzWCAX6rpOx
05Rh+/FlBZ/UxQl5U2wbJfI81QioI1luiWETkRwgZq/Be/tVKXrFW/3bexllB9QV
0yqRYI3sJuQBhZsoSiYidQMTk/Kd+/TRV3Wtip4EwXOnkU2mcIUKd6gJqH/qUkHj
7zVdIomC7j2k+71CAYFjn7Ryo0uekVliLK27Q4RSqMsBW830K6fjzsuDuCag04oG
BIEAIGn0Xo5egrANV4XZ78WceDWIU0Dunt+2EuYDNpart8XXEk5oWTdPTgUhA57S
EC40uOuejNXJsJR75h8sMck95wvfhGi/i6lJZDnp4j/CMmj2MKlr1nIh5cI1yszd
hSE42LIUdkLub0X64dd8daTCVA3svLDuRQGOqK1nGSbt6QmoV3iPlfuG7RhOzb3Z
HDvYTXdBDmr9kGl1BPFVaA1LtuDyIawzvKIixgUihZaLfpzFJ4IHpM0V/9Di6umb
fK/XTHTHQmfpiXffXADkpnbS8sLa/jIrBMSWgy+JfRZCUxCEqKBHJ8prQZ0/RC++
e2c6k8qNEgwhCs6wp1lRRaR2VY8hE5KEfitu7xcOOsh5ln5PF+0QYSyjTA0Ywl/K
yaLdnVBt79pzQUxOChHvPoQ8g5UraLBpY1F1VSovquq2A9wxiWSzUy5F0tc1DMWm
TiZSNaNpZuhY3q3Gw76/7wT1jQn41oKbTAFiKNdqSPpVjGmXfkCp2dcRtUQVKBu8
bRqCwcrq87xwWMLYq2E4YmpkkN2YdEenuSDej07/gG33uKq/URI8dRVdm2q7taq5
eeinvpuCCKa16pvE3CUhYzLqxalt8CUB6zw32eGnb1WayP5JCL3cLoP73bX0TQeV
r4basZS4xb2e8v3vkGwDNmWk33OWBwG6X/WuwHaajldqpUCdElPSerI5srhb/cie
P1CKOYzmeTXAH7x1lrVETIFAlprZaRUqFVT8ThQL1c05GR19b1/x1HHGFrwlKe0O
4b+4gAZHGxCpP9kmRSyWxCjE1Sj0KSkmSguBxEEqEzA+uheVV7pQxbKDIvEcoqgi
iZ0gBpFbPf1JNntJ4zlkS0r7FYxRKVRbd/nN1M5Ho0f7pzP+Q7Jv5U8+xQCy6OmV
lnTg5JTmlt4vcpoLBsDRk5vDuWRKSf6hKWPV5oUqhUJcTWz9F2Tz2ZVEDetypuln
2GjZ83z1wMtLFLG5+HQiw+Klk6T11CkN9fub4NZMiBIvf/fyHakOfuWlan3bsmTX
xzGKYC4c6nPtvjLlIF/hexZTnINStIQCW4L/J6Atqw+0xy6wCOFAX9YZjHunzCQe
OjMRWwlf7unKdPh4iWSj5ULCLqJSkM7RmDdn29KplXtv8d8qnzK0uenmbWFsuURM
fkryDmR3dY3E9tRTfO8vfRblg9UQEcXOzGOmgGz9Gtj3DwJtN7enskqxzr2eviqB
3jlCOktA0E+4M1ykJY35NAQwWHRnO9zC+zH17IfHiD/GZSbp9tuNjbbDpbtkB5de
1+RUv75jP+nAfR9YK40CbGxv1QyEmbbfaCsbVwn+YXYxscJjzZSSldUdllcR0hRF
3Kp0b2Wq7yOExwBNgSZuVk7ayRPB+SccYowc37pzdQvpO1v3v1XMi48YrEI4GYoq
DpF+5YrOxG+0vCLIETYCCdI1j9arLXRmOPxD386pYKY9iC8FmB1d8idmou45CEF6
z3JIYE+0+XlQug6k6aOtadDIFZnBAYsfBKMyPJvq9ydmW3lW6zsN1JoyCp0GlPFh
YguZsE3Q81ohUmKNMzvz+hEbyqd9ZVv/x7sPrWG7rj7qWr+sWP/cLV/8g26Rvxk+
+G8h6wN+AYxUU/iI79TFXsiw9kSGVPRR/XAszHYP9wQV11QVbjetfufQJvFuPnSl
8qQsJFUROymAEH7pSJ6VK7RbaGdBHC8ZF0YrC2XlwAm+N1gYT36tDrEGteG4WjYD
bjHX772xWa/nfzJPiVNaPMM9acCocTu89bo4Zw+B0BRBQVXSzqEik0DXl6Y8xVg5
ciAZnMbzjAElgeYdWrHgQVtItqdMHkBQHf5VZPg/iEz6NmWkJqdnmLWVjPxKcVky
erMwRRKA6FFtbXPcOyOVQKPlxi0F2nyMfbngqPm4pqG6Jt9tBU26haH5yGVsUJVJ
TlVPjgUzqnx0rADmm7/D6VoHkQuRHKpYgqyu2KTmiGkBa0TNjbIuTIXskzqcb89w
jGHv+Kl36KQteFAzLoKtPyDgCXQZhdQbZjeES8xzGvcZHHu9o3N2fVo3JJXe9J7n
2V+m5G9N8NzSTaK0c4uSSb2eDyu2Z/MYjGdeuKM4floIrCIWuOQlOK8xgz7wMUBu
Xd/JUu5Bdau/iLV8kZDAXpe28qrK44yyETPUBG0/214AzBUEbz1P/KxG0DKKPX15
M2SEFq1pqope+Eo3H11+vecz10DxUrF5Gh/HrfAwUIlP+9942Wr3siShZlW/NZYu
SAAFIPMWyFB8oJp+nz4Vd1FLjRNC4FKkss+7l5jA0ias7LVnvvWUDM6GQk4fioon
7lK/rbK5aZO41C6zM2rGjBxs98WBZ4cGa3jOGpdUJN8F/8RGAunebNsdzqr07YfM
H/gR+89lfOlvaA3ik9E+EmPyjSGY2rWBRKftvt5bfijtNisfbQ2sCHnzrHh+BWBv
dqBa6mT56HPUofblj1kLN+M7LWzGB8z/t2HGcM35CfonMLz40S+nowYO5+RqEVHq
cdSNSO4aUXf+lgJIRstZ1VJVgiFCADPKbh1GLLbF8kEp/Gk17NuyMPcRwEhJwZpH
y8tdj5A6To2a7CSjrbAZ40Szrq73+etKx1DwxK2jxAFqA0GTiePje7ROjLJDZL//
KA7IA652bl90jJy+Gb/YZT/DuWLuuA7q/1E4Ua4GMpAV2yRoUA67H4rQQ2PNyrNI
QK7Qa2gqO3zJOZBvPLoCzDY3RtZqFni+d59/x5YOgQTJLk0cQ60xkbNppVrlrVJp
8t9PYbR937rHiGqqnYZzL7U+NRe4VXs6yQ0cz4DJZih/VkC9uPyNTR/AGLvJBOnN
MkbIYnzy1Yea48OI1/tzyqrv8bJApSaMVCWKmZ9ciah223spGcgmH39IPwdxFhPf
HKQC/ZAnk2xSfYh/csdIo59AdKyB2bwhm3yL/NI+DjBKsljNZYBy+KQyT2nVDGM9
qgUc2Wd6tQNvBfHyGOsAmPkgg0eT9rvpjzSPMmyePOUyr8DTtOiKENCTrLAlBx96
/kq4JlPFy0lME6Q8glSZrMnCOEhxOyNIH9Qn4/KuWo7ZhwxmvyJI0jgJLnjTjudO
VteDRsm1yel3YOSs50SLXObcLM9c3xW++LFrwQqcx0e+9QNSB8707wnR3d7aPP/j
wXvlNVxiiYagWDHsXG0tv/2tlza/li7nEbQGxNiavqPOjYLjTsgNRONB3XFT6fIb
E8GQG81aypaBh2sF1tFoC+92GoDQ1T2ZQEwkw+26hxT1Shp8XEfy1w8Jjy5ABi57
tbMna9gtVDoFke+j+qny7rAUOgMIscBm50m736lw4emCDMjNxnXMm1gbLPm+JoTQ
8g8XBTXOUF9zbBxWvKkqobWfnRvAC2VLRE8uxa0BJNyLHs5+h7PfY7LoT6RqZCV1
zml3Nf5cbCzNk5AIydZ3BjtcYzHAksCWs7+DGRaH2y8yUkjnREIfp0AscEy76/Uv
Bl/SlFvFCkGQmcGn8zJf+2IedmaoMj/XePOroWnhbi38UQwO1KCfur4grPQ5Z/+F
IsmTGjOXjSqcw6Z+qT8nCRcMYZGUEjGAIYAmSNK2Dif/l+CRm2QqjanV/vwE9iF7
8+31rwmoPYsbt8pIoS4yaoOeVHm5wRcUeyFlr8hol5FyoR3AstIy2XSsWbAqCJNY
z4ru0WyiRs9vfaEjOOhju3Gqnvqd3s5PC5WGXHyxphZ+LlDdzo7pdVAfly8MsmDz
Sr/Mg/2LFZsGq+OQziiaDBGIF6V9uKRz45+QB1iBkafUr3OGTSfpGFO6Na+47cC+
Z3TgTTAFkd6Td2bkgRDxe7GtZxXlnaYQN+/6ZWs0hkqxOatS7v/VoKpfyVcr7gng
FEX0jX7WcgmFBmWQToK0BBsnTc7GTTyhWLD07XtS27LRMHv765nCC8F2eHMNI35e
WTs/JMZYQjhhRjAPgr3xlzROquMbIS9zPTstg0CRqCAdA72r49Cks1t1zrYoqXYr
+JKw8EjIpSIx/V4wG08GmaADntjHnt+ceLWc8A7fyT2M7LxBvHo2uzcirplU7i2c
UhMBCMKzDoleaeBt2RcknmY0x1mZKr0HRH78b6kcBqVOLVsQ9lS8YvZv5Tn15ib8
f+mQ4+WIw/JSYCIn+QmObgQX36e8ZtSkc+dnpGQ8Mb+tbIZhKKpzTtQg2ieadmp5
BNqPwuBmHFFU/9kTnL93531z2FFTkKm88C/ThjAG9RJboXOIsxoyy6vOcc17gY+v
UWwW8kZSkay3UU+7qfCDvtcZUFiZZSxpYh7wsBusrFeltqaJuMLjcsRyK1BbN6km
Cx+03QRyjl+wu84WAbw+r5NEecByoleMheQQFUQ3S2wryuhIe5n80JXmwsr7tB2n
Cc/qKgW0wFOWHfE0UWd9KWWnFR+1KUETrcr1NHUCQ1xbpE5YjM6lWZx9N0GjMcma
KfvUkgEq8xvCDSh3TRhryIbBh1X22/om1TJ4UUeOUcnp7lAK9Xrpo5gsOdt3rmqU
z2CcKFzEvnk5EihAGfkqjx5xErvW8ex0REclCyfhnxqRd+KLU5+oEQNLWcDk1wY9
XbZpc/UbYXRmYUPo1YdILZl0lPEwuYOXpI/WoLVqK3gV84xjupkUXVbNCjSp2SO0
3YXmT+1VttdoPJArCzRrmAOMsKQyr8pNF6ikyLMQpQ1icaIij+dHeAfmYJxXeegY
dc2EXlRTH4etf245c7I9cI9QnRtFQsfOImOKLFKvIaGLIfWkk+L0rBnVjPGjkVDz
dyLF9KizDrg8r6J+9wXpHPClBSUX2qTz6S8tBGJ2RO1E7YQAlhvO1QTmeb0LbpSK
YkecwyT7B42XKJ//LJ7d1jWYRJS2d7o31t3Dv7B367vbkhTIm39TNsTFciCWi0Em
Tq8hC8RELcZbviHsJzmHwhQ6W0yD/D8JpmcdpYhGDRh9+qUGP3IxtOlLKA/2+msZ
Hcsg35CT6D76apiFV0956bgXL4XGUiC9MsmZJmJL1hWrs3t6363F+4NZfdGxMkEJ
XI1SCgmryHJiCfeZtVUf1Bc+u2x//HDOPbf0CHrUyaGo2E0A3ztJJ8ssJv2beYGF
9v1q04TnYe7rYpE0eJdGPsYDNv+2Xzpmhi+7wwS3K7HJFey+Q7MRYBawO8uDSTUk
nncz+v0TsaApxOSfuqqAshMpdbbjNQ64flTWnvIjS7epBy5FsF7/NTfKEObMrdF/
O8sjei/0PfORpG1zAJGp59aTOjJbIU4/HnlK4JagGl7SIU79gilRzAB8g1aJUTO5
yWn+y7l/XRiKYpXdaRVUJZHKIU+bs3mAwec956T3N1dRkF0YzSV9bBk8xqXRMkHf
+BR3b+3RfVZad74ZeoS/jyIhLAptb8AfLQBMb93MQGElVLl8wbW4QdPppbwi1bSS
B86vaQ3JwfgdO3sKevVsld/WqOv1rAGHWSg8uxNMzD5j3qx9Gatry/Sl7dVpxlCH
WdUbXipLkJtbGthHHTlLP055h48JShHiRpz4wmfRQUBO/ggWHl0rrklaZVLJmsaZ
kt/TKM2+clk9c8hxCSVlkeyENpK1V2yJtk9zXJc7XmC3fpHu1EHLUT/RfIar8cEe
KG18Y1rVisMOu5Ha7CM+c7MbTJ0lz1tO5VhodxwvIuEs5VPSrxUrW/2Yh7LS1fe1
0UTpRUrrVNc4X5ixy1brlxdD/G7jOjb6qeb0epqbzt3h5YpCXww8XkMRb4tTeIxK
VhNLKkkExaqcT1ORCg0TxAr93EiMS2/Ih9MBbSeO2K8AH0Z4l+1niqnDcDiW+L0Q
4Tw9LzlN152ZOKppWel/GnGGIcGqUhRvIHmDqPoDDb8lg7sLCvFzdmouS0pc88Yo
31TJ3jdwYb5rGZFHGTfLfpKaoZSqsxiKl0ZZ9fLthD9+jgMYjpNPMM1YtfzmPTF2
0NuCLJW9dJxD9FNkrzTtfAgpSwXDq99QQsMFYHhXZZ0MzLgJeZHV/p5GePIYNXGT
xYUYtKuG8/aIp62mqjzUImZvlClLELW5tRfyN3ujfrsgFZMpEmLQT1AFEiJvT6as
8HcF4KP1WLITaP8xqlHVxK2LkerERPt4CGyAO5Anx70caRmcbk8LZz7nyupE9uSM
japTtRspWC+bXtaQshd4wZpnajhwDymytG2vFH7rulh6vB3C34J2adpXPyD1df9L
U5B1WOi/fol0pilwWARRFVrEm7IgeifQeEy909Q8Gfd44/safDvBsGe2mOEs50rj
m+gqyf5jn1kAvqNn7C8LbHrnrPI0GckIAMpLrj3PEQ8Rrf1tubnuVtEC7XfgrWDc
uaMiWsiPL+Mou59/bh8RbQXP4iFn9E1Ldk01aWffFQc0OJcPnTtaN6ZVjAJU7sDs
ZhoUvcLKbMQcHBqda2YrRmWVVn01UNICczQsGV/yoPmCGFxvU1SRdk9O7N8g2OyO
CCg+U11X/bPxq2HL3IA+O3FRTiOkJIpN8Y91iPeY8HdleuKUMfd6bUYiv+xnSFPe
mP8o12V2AvxC4rr3pqlI1c5q21EKR7sU7IqiXrabDda0YvRTQkXiO5pjfEFAfBcT
qtjoQ/OoBe3wUArGkaMe36H0PpTXINjzLLxSas5wT1iDcqjZ2pJUG/lUeRS4I2Sg
cu/+DPky2tpNxlaYcsDZibx6WLg8sv6ZGkpgdaNv6ArlK3OpLqdbNcklV3la57sC
gmG4VRITsIcAZy9SC8kmHIEyaFomQpUbWN1b6DjD3+tRbtBdlUn7qJVEMGobMT5Y
Ad9Cy54SkwU2Ar8rVpJAvzSUNFm7gMVidGOq+lg02JkrK/wIy6OzReNIlBLTXGO1
wWM2hUYqRVsJmaeQt3CiYimCXtDbrvpj8zFC1nxG+TGF/lW7KV8IqIDq93QspH6o
/Y7W/58EWopsGQiI9+w656hEBhRMmlG5/cHh7MJ1uKKaEe9bz7SVcYMyegqce2YO
FaAmIqechZ1foKoKJPSIexev8MXZEN0jCxxMcTeFdIUKWm/bWD8F3VUaPitLiCMs
Obv3aYXJ4HJuea6o+E7f2dW+HkD6siOK4guH0ABgqejwI+eSIJrL5NCTudY2hiu2
eO5iIA975x+/hr5OhUAzCFUUdU/tK8o5CSVcJOAN713jqusYuaQT76rcyaKat3Hw
Sc9ZKVRKefGSctjEgT4qRNNgxy/4Se0lNmQNDUBgSAWa0yvktmstUdj6qlIZbv7G
gf1c8v30Nxp+DFlBs6nnuSamyMLAhXXoSC5cnUz8pWlIAW69/yJuUNq9Dv7KShuo
K9JRF7uJddmoQEN1K1t3EzNznpk1mvjizvjGBusp3nk6MBeHjN55KvIizn0UtsoC
5/AvJAVuexpBPjqFCGlI/xbRBF0srlX+mC0R4faU8co8p2gdfibZ5Sr7jyv05Gci
JjTsVRgfK86olg5xLlZ5T5nBeOKRyYA5trFiU0HCWxmSLgS4iZcHdFZ7WuScobHJ
D0iVpOzFxM0EJs+JU8oILxV/JAWdWoghm1WfB8XSCWALkB+ysW30IND7OHx+TGqs
j9m3t/jOnw3qmFj9T8m/Js6yKfuHDt/JuSjCrTnfxZWDv/LpPXHy/o9o2AX5+fay
zyE8z7aJy8cZsHmPKQilg34vO7n+saOL4C+1fyJBC0ArGtCH5Fi3oi5oQD+Oxeh0
GXmuH+Ixh90Z6moWU40qFyL71t7RAOXkQe/ownlAYIuUTOA37eTnbNBHUuuN+ZNb
vqyJcRRqr2yRYJzFYMDrQLF2zLtq0+AB/bxfpDGByMqZaL4CrwlZJwZzgjhQxbyP
H3/UNvFTlMD0yzVScQmnPjn3JcC1crT6br9otZXOjxXvH19oEdi8zQmddQ92KvdD
LSkq8ziWngEET4cmsAPTdYjewS03zDjWcpqUv7Nr4Ip9ndl/NUTS4RremxlCj3mv
76Yn8XCZpZZMSUQLtpSIxcOefGlZFZodWHnz9E3q578LleIc1+NNwPqMdB66zaES
IMltGHZI4Kr/Ik9w8LeKPJmEaJMspaXNuIsRWe0kr3DD2uCi55teX5sW4Z/Q5rGG
soM2t+jMTd8pC+ncp8vXqKJgjsXlwvNUDyvK0GIIVOaYrpzZ4A1MUZ/hyJcwe05y
nFEGu1MgyhH2AfgfLe3/sauVr7A4O1N7ulyQWu3wqpA2nEkVghUDV3sfTtdf70u5
e5icq99tzskmDkVcYFCt5YGCY9XndjMRqzehDe4/31okTE276ByDGbn/YHx5625S
J5M9wjwNlS4LP/HuE8EW3DNr5sfGWDtBpRzB8EFohrAybQaujdeab+fq/wUV3abk
h3Nn7pcvAtl5jyBKQN01S2BFNJPKQV1sl3hv1mXi+3s6x4X4xolE+OELQwAGjjhy
+MDgXQulo0cxL2B2byxx0HE3U8SC95mSimMZDAakw4nfvZZ0xmqWrDf+6Eu4DHJf
L/3w0DilcXuK2ihpCg1TVuPW4c4IBdsNy/ICgzfobQU2jug/X3rni+BeT6u+8UJT
z4ejwAsvD/fezsqgC3Vfdg57myA95JxpTmspF1dcwE+kvYx4ocwiU5hnCFZWu9PE
H8NYNMBOmtGYjHQW3OTuVlyihBZgMfIEHgDQHJjicxm9BkgHlQkV7r9+mGOjka5x
c6N2VfSdz7cIgoRE/lOdLf8D7bRawZsSTa9zZZzfJ/5hnYC5ph91pd3Z4DpPsuqu
bAFBQlpj8QIy79ArMOWmDuK7UIn0OTBqDMJ6lJB72CVDfNtaqZv+ZJMghgYIJh3/
EqzJJJ0PhLiSEx2w8+0TGzSJIracB8C/D0loEXeqU/d+skEESXvfiM7uaFhBjxA4
P0qht74XD23MGyrwx1TpTeIji+4vyk9peS9wjY5bHEdJAJER6yewzziyuqUsb2pO
W+A6bm4Mpl7BcIReGB5+6Mu8LPddb96z+/M6WLDj0WeKfAm0tzdrgjsBvw3PGIuT
XHbzXvviYSY8oaWOLe53ujc3bw9T2bB1XmLJxuxjxn6+vBPZtQIQd3R//3nc5yCM
E71e7PPDxa8p6ecIKskCG4gOgH/OvJT10LJgUnfT4/PkfAFUV1NXK6VI0/DBzaCg
9YPkvzD1UMerz0zdFitH0saTbX35CEfH+/94Q5B3dbpeYWLi4Y45VFj+rohQwIzy
8/dSSFex/TlEGWI0HVQMtXUCJ651XkePCv5JZHZEZUBHbn1cpgkZ1aQRUNLKXMbE
WQr00mfiHep/KnaMgAgbvtlwIDK9coq0gG+4gRl74p/I6ErAJPnLEiGovhNh20WV
Xa39FXp4ws74aOn+noYuC7z3dOtxI6WRKXqhkrnqRyMQZqd/KOEysZzbS0G9lh9R
kaCgkDVyHin6B/66ds632TQC3mgC7Ln1bwr7aYQgw3mtDyVPdnetX/OVMma00n4e
CCRHm/nlIQ0u3H+NB5khfyfbRFVu+JqIatW/e9ERkEpeITJiIav7dLXJIh4tRg82
saJhUbWpG+PVnho/zTLDRaW64Rx8gzvZKdI+rY7J/ao5VOD3Go+OhL+3GQMqbZUC
uxsjN3q7vFvpIbqdhPPF2sGALd/jr9Tod0TS/ENtpKh9kOQS1Y0LoWylAtCm9vqe
uGylIk0l6+7X5s0tcVO+3PQavbujPKqW85qN2V2mUiHEbu5l9JXxSK2A521urbyU
kdLnVAD/tWdLqLBckPOue+WQTC3ax0q+WrAP5ceEP4blTEv3Y7plLlQHLFiKLcH1
hD4MGj1fUsHqEhEtFn5K6w0sEZU6IQ49FC4CvfA+G3SdI1nHuG2PYYH5oxEp9LqC
zWdBbYDG8Vtdfzsczt4DJVBf/17DKJnVJjz0DK6ozCsi7Ys1EhAV+M0abW2h951J
8/XzH1xwG82I53tzD6HNLDRvqdBEkkE2r/IAB+s1SOz+njniZgoWr2q4rR8nujm0
8T/CTUc2p+prZUo0M+sTXQYM3N2D+mvcofPBm+O2BcLO7ibaZn+FXlOHNjKsatIl
uQVpny3ot7gmXSFBzpBuWLnw+uiwRPxaARcA+mVmSpjzd4HBZBSXAs6w6OY+4Aki
8T7iH+YzmuUW/jUaAHbLeZscLEk1hNFhxifwrtAK5JOZM+1LDJijY00uFfEJxZNr
GVcw1IGdy3hzrW2MuDUgjWzSI8GWGvyc8kAfxNTKie6brHiHEKhMOvR5AGX7pdfb
hcpDuM7RhbC+d5WGDM+dQh5L8+XQneLwyofrnEFpTqBU3nVswnNyDy30C68CcaM9
FiYdvP/ATJOscV4hHWuxZyBEREtYw+ISkTJP3W60AagHEmCdPwGzYdhkg3PSzhjQ
Fx18rU8nNlM5lujcqTemRc67hG7KqvIXoYqhvvbkTiZbjB0NuknDB+03iLhcXLEG
SaivyAZxCaXL5j8a5bXb3Qd/9/nRrlvNRQbH1IAHmwlOETKyU5Dif4dbe4BluSHf
xVZF+dso16oWbH0B8cLMdufq07wl2+DJTA6dFGPVxPkZCTMiMm+Teatio+pNfG1V
IOnaT6qkJBQAl9kLnJ/9jd3FYTEqlRzeXVL8Y9MNxxfM2ktK0YqOLxyT47hXgPXD
WM4+8xiOZaphKwTmJ+//2p0xiP/f1hDcv40wkDglUJR61Ou1DAwAmfzSsysWMQIB
wiM9xauE30I7AYPfeKlGmnm+hlRpvx5bgwa2HVzzLHNcgF++rWOONf7OFzlwPni6
xLDhddmzFHRzu2A8ShYe+JM7ArxIsmBnv9A23RX+gsMU6nUAQuGn87KSFWTVp140
IuwHjrjySyUoKg3JJmmauYhKgNkDIXCLPDifuRdrfeh5wXbQR0IgzGJmPhYLHBuC
ojPSIJ+NTQtX6RKN694lBn4EKHaVMyAfj8Ejya1DJF/Xv/yT8k+VP6tiq/rm+Dxl
SKpggDiYkLyvYnmi5wFlcv7s8OQryXd5YepklkwCmwjCL34odc2+2x4IEMOhfXij
o5DmFyRsIb9wH/Vby6MiwYhb8jOpVdD+nubY8+t9yUpPToA8aGFCSzCDWE+Z+KEi
ra7v/PPwzEabDUJSWtA4B6/d/LZfdZJns0RGUy+qw/6xEZm54mO1dxyJ0eTmq6Pr
hQJfX7ZJzpn+2baj2qopESg4Kt84gn7fl5Y1ysggXo/XdmUkvjDVvmfc4BlyOWWQ
oQ6NJtX7wH1I/ZoiOsXCGbfltlCrR5EJUO+YWXR9CH4V9iPULUAUyeeZsefZc2nW
J4c73ANznSa2l2tID+HVsChNQB0HdFfvKTfzmd28i7SgJSAi1PNOjuBb1qeckGYU
I5WzvdZb474lJAEG9tP0vaLTNCEIfk+tsMaPFcaJhtZkOgSbhnE7SQacTTULf83p
9i7+UMBxnLexaCMVTbYtKfiN2LyJ9XDkYmGlA8PfgJjD0JvaOu8NzGkv6H4tv5qE
jV/oYnb6R4GARqggTnBCTbbGfvrpK1JZGfQPtj9io5H7xyK1Ol7OKjhV+q8kuZv0
JxfUxnCauGJyHNoKNTca3kUJzBnJ3HgaqPDYxIYDoqIWjYFQZUNdz/o7YbgW8cht
zemGNI/VtCTL74x8crwc9I1z6vZd0B8D1fLYURZI3Az4kpOYiPFTTwK8G76Skqpw
llaPs/Z1orC0O06vMwAifX0CMqfuuQSNMSH+mxdkeUgpypwau/CjDihM8f6nGs1e
lma3MkBL+pXxqWl4j89EEGkbZ3SZAshWVaohayQUB9R2i5Z+G8suBaqfHC84kZFr
th63b/9gdi7X6RaJqWZ5m5MHaOm7BDUpqDNe6/mDVv2tGY6/1SFfO6lX0yZApBQv
Zz8or5t1eRuzA7k/6LDfbQuY94AtXU6ZT+yY/lDiL/XvBQYKHodFkBNJKNkij2EW
O0YsqJny4H2J6KQwpZyGL1NdwGqw3iDguM86GzcpuOO0e1mo+hW/QwRbhIMSjN4C
n1NQyaixlDXbqsiH2qJCFRvtwkWIZGkUpMtl8xII07UeKFA33qDbF5XMtJMjMBJD
8g+wo3s1AEbQ85f7Z1IT4DT2QpBYvkITz5X5dYXLGO59iaf2HSrZXiBjeKFT4D98
D/41J/Tnh4s+VqRTtFflHkMgRocOlDvoYTGU8ni4Tm7jy9sQ3zb/rwUyf9IfMhkn
TVIMgsHL5ENshdmdfhN9BcrSHhtPt0ZO7bTpIsv1+D37AwVwzWlV0mgwnXbEBYjF
XKXlHBdVGkBugNpUE9hfSZWNbipq0XwPC86mjjfCzlSF5zQRzWZu4zZM4daW6JsO
0Ba1DH8AN6RgP1FjyIQc39tIzYiU8EgW1s6B6+nyOm9JErDc8Fo5tY19+VgXvHUi
vP2wl95ipdSUqKaDVe7fLCbiv8mR7I5uOp2ykLAfVg+ZvLpdAAAAMih1qQ4MFTqx
h9L+X/xOabm6Qz227NstFmK3CWXAe1CB5wyEtsEJlJ/BnpIZJxfPgNNPsQ1O4hr7
/3KDbmPiltf+NHbowGJNADkrfj63RUSqT+7axzy4+Yx350a0xZtm5X4HmC2E+6fJ
VVCsCkhXCZhXHygLmxB6p26XwTgk+M0Gzd9YjF8WLlZcOb7ftCU2PIXCOUGLimsz
H5ri8cU/C8h9qqpxtaWOfgKs36uEVIfkRsA8HXPCJsDBJtc3iGpOHR0/qWiGfpz6
m05x6+zZFSvRkkfWNJPWT8IE8qFHW0IkKd6UHdUcZscErIGMYGjrGVSwtcI9Cvll
DQL+v8OpLliZeU1dnJkZ9je4aq6pvLOslw1Xw9o8TsI8zszJJra/izZU8iswO659
BZ/z8LUg1lHZ4zhU8cxpqy66WOae+VylCDCoSTNdMfzpeIAyOV1oDvyz25XZh+HR
MY16slxmPUOJ/PlGfV9Iout0gKXG3o2Z1pNfYlAprdv8LB4BwJtkyLWFwhNNpQsg
byp3AVk/0KwYjgWi374N3hBUOfbNo2BnQPuSKWm/nwUnHu0gRd4nX6NZKTPOMS7w
Zdx9weU4945BwMU8TASC5jl4YOjbpGqdr9jaRtQSrPpINWgXskRcxj0veWtcl0TV
UafN+EWKsgVAG12UZPmXuq0OkFkpZUtAciSlChuv22hWQC9shYWmQxxSLdQdvBoI
Qw6yEurxxa8HnHmQy16yZQtZnWxBX35HowX5MJdbJUIfK8heA0HdJf0UIaxWixD5
KuUEqaBhlMVc83rLzDf17xf+6hsOWfK3I/fRzPSwbRYNvCuMyg8Iw6kMNFBuXVy9
T1hm3Xroyc5CljTmAuG7MAxoQwOu49LVFCLlL6YOlm2YPSt8YJ2nORVOs8ZvtjpX
j7EYUKdHcQXmNB17McYFK34EjF/U0Km3LRa+qDDNTbVshGA3lAQCWJD0mSwllS6O
BQIU85zJgbYzcxFDXk+J7prSR4wV/7CFl66MAVrgTRjI05eDBic9z2aaRMqQbwi+
8DvbCNNxpFPLoQ67n5itHPlb2pr+2vfb31v3irjTtP3BTbDQNqzhTY2gdcXDIzaA
682N+QRKELhF+mXkqIBf1hKTPaAE5D94vDNEdQ/ucCz7iNWBQFFOEpZh6OPx/42S
i+FBb4tiRZAmy4mNstfqZXL1xvpOF/BeVtnifMpbcrFa3yc2OmOLJHynvEuDGMER
doXvFUpYcWZCo4yL2eWDckovxKBJEgx91q6XISZSEEcRqCeZwKZgUCWAbnOMac5c
hKNDRcYq0GrKFHKpsVZRu/7+k1WHeUEHxJLXsa5L2DbeFFBMVb0OQQ0s9b2KTZ6R
ncKKOM+ceRf5vlscw8J2KMDVrdR8GnlriJQC4iYM+gKIQTaREe800o1DPGE9+iHq
wt05lSj2JzjwvdtlQ/RwNV0/GTMDRv8gVySqDUM0SrDXn6eIb8Uhp4pwtiMdhqYO
F7V5g/wQQjX0dzkonvC4HMkVa1UnKo7cl43JZIA0KRy6YtlaFAQa45bMsKwHJ2op
6Q2UjpyKnncIrgOygmuN4ip/4diulfbJBLP/2vVc0iZJQkZFQTShOC9Lt+O21ax4
Yo6vn/wiyyy5KtzznJi+yUeRVhrLd0m3asNyAPizDpacSZ56ybWYDThBL41F2QKB
l4+J7xBO2FWO8nhTcOSuieIYgrV+fNQu3JLG0lR9odlnwq+i6IfZ39Bw7yhBjtRS
IlnnNZx3kEwRYZH+WGovF0lo5USdxR4MbCSXn0FfBQhDtRZi1VbxkJuSjLnO+Doc
VX9t1aUo3z/qBBl6+uaL6GBS9mJV8OnQYkHb4uwHI7j8vQakn9xvx/wmCppjohqk
eKdnFdFaWlV1UW7jqmS4BpboFsvsLOarktUtY5KULsOgMRwZ0vjfx9NTAyKhQkTi
LkxgGKuxtbsWtGoj/i82tdY1yV+4LT64+Z6bAJXQLOSTNNdZ9D4GOzI53BV3nO6e
Ls+NNbhgRjKq+uEbhe2i//vhu+bBxLtASJ0rvOFjPosvjHc3rNvBeweHMHQ7N2QR
gEfITLM3pK1gVmhI3BTQDRL/OURZJh07rSbclkro5pYAbT7AFoAhlXlt2Jli+AiP
iYLdCn+dUAMPwPDCLJBJuKeTf1CQbL5thPEllk/TuldYe+GFTJUXx6mB0kLugZt5
uP03Z6YvitrKVy5lE0NJKS9VVm4QI8Ma7fglpRagRQAhWbbRbLoBbgR2UyDb/dfc
dLhcjHFz866tfwFLKUvudIkiwEg8VY7iK/8wmmowlMsYQURj6l/2Uk2UyMrUqTpc
tywIGZz+MmvZayM+lrLixDNy0PJzxQPZZtP3I1tMUr4SxF8lLIkbuHqS9z6mWQJY
GdBHGKBTtpO73LNkuqFaS0fh7yVRoeAOo74bNNiVvVMk95pKiXSEZzjv1iTAewMt
IaCUKJ9f4nogZrhh3ARnaGR0nqQfNjl2miS945lJ54B2xDjPZjx68zvOOQSQbN/A
4Foie9k+UkGPnpYrZmNvzDgMBp3W3Lbcy6EO0hwctOGUy38FodFPg50Rf38kS9CS
dhndlPg7VwFSMGs1RehEYtVK7cqryGzKHYvDJV7qxLDhqLURe793x1CFbq4uL5KM
Oovnw3s1ZydfILdOm/sKUiDaVu4Jo11wzuH+Dvu70a+sCShkB6xBJQipXBje7ekj
mYHeostVI1INnOeFVkn2SYHPahHLHG4+96Atcp6pTR2jQJVaCrI3YdPFoozfKcV0
cZOFZix+C+YL3DbbrhdW+2ILWvskKMLcLQFCyGpR6U4CRV94dE9IpykuydnRjMSQ
kEbiDKGzoJ9HSq04pl8/nopu/3DMYx49r0pladwGd3lZYcVfEvGK8swws/CkEof3
nVNQBkESTmSe6Y03cbC781mpq2w0U7nehoa2vhzfvHiB4Gidr/WMoHa78A10lyQW
BnMYc1lGwcnEIBtt+4Tmn8ByQoWomoaZYRNuigot5MZLyAToUpA5u3mheMKgC4oM
iCnb8rrCGT6eHXYwe98XVlzrgcJmwQifryWwmq50OUYpO8K9adCWjN4tCKtTEBZE
BnkayIFlA5aj8BMn2uTEtg6TjNtK9Zl4t7G4tfo6KKdTCbMZrM5MSPS8kXfJU8qo
/krHfDXeHXXiRdzCJVRZIfMuSFZuxFTVvk7bAorXFABDp6I3QAOKyqU48XnkiBf0
TVIZeggWIsc3iQxdZFYpkIbEQv8fU3UOPOGryG5l5Ln23uN/8r5ySxiBH1OV7Zgh
X/F+jTrRC9CTD96wBuvfNSA7+qYgkEMcTaX6bQE5wkT+bN+olSvOh6DbP0p6M66y
VYphXLvb1+IquT+VXBFMcoqUATnUNCo1BPkiGTfh+sr2jNO7DFXJe5HXKFRYgZak
2jubnd8QXaZCylXK76de96Mo9VnLmBnedObV1rc/j7kcK6FLzH+7WSF55tMRJ2/k
XnkvVhIPSGh1KK682Am3o9E5tQrlxZJvYrrei48RpWIwUcQQxfkM/tsR5Ve6SNBs
ZjqnDOZzW2GhlTqHxtx4T9qMxrfbzoZsUIQu+4e0gwePRN6ys1ndKnpNHXuKylnt
6ifMhbRop6OSrltc9zVmlfsI7eBQ4MV9CLDhqdWkPVKsEl0O8B+wxd8oM850V5XT
cFT/Cue8JZ68w/3LkpoNIVAaRFiy5HDMQ75YUvmMzQSgyQz2kyd6kE2MEb/IkhEo
PSw0ybRP9d9VPfIuUl/2SzkvT1IgpKQPzM2jV7/D3zSZ5/ThKbvpBoSrgAoeVYh/
f+DFRPXz9aO14a28HQuQI7uPhrwdTcwU1wx5llYJMJBXS3NXIdatOKDpkc+zrfYL
BPIduIE+InHiCn0iYYsmmpX92g+/PFqr88PS/lnP2KjcWAoaLXUvoC0o0aoyjzNy
C4jjZ9uG7feYp8KRvpBf2wvpwa/VOmYbFwwBsEuDnNPQohMw++CKzZLbYGvp3/MQ
mZxkCL7IPqoANuPKCGB3fwBw90QpHYbDQr4Z2E873nbWYkO/z1xPBS1ZOzhC2y7S
hwHWX5O3xWvMISyRQ12N40LqRfIhpK1lyJdVd3n8IFMejYYpu9YQ90HgJpKAzm9J
v0Q9aQirS5qDPVdznD72QEw7Y6CQTYEM38KvNmhAPUEhkopm4Vb1lYRVq3OT000q
omWG6yTkHI1WWV1jtEzBrXP91QlweWNKxCmnyjS/r3K0S6WA6i5J/WNJbGv9gASj
FVUggSvkpEPZq/5Z9IwkD8x/tr/xbtzr2qitFCBvNYSRzSgkXnaIKiwX7dZelues
7r/C5weB+Lwyxiajlv2wsMIxLIDsU/18ABcyxa1VQmwnIGhocLS1oqOTLZKohhs9
fMS/IeSzUR2dkaJEkDeZ5Xf9cNDMx5z9KNrzUqe5YV3zxMKlqA8SdBoG8sy+EpJ2
MLkz1SzjuwR0X3aPEr7ZtQgovvES7wFtqpno6CxPOKAnkEx40iuMCCI4NiyaTuhX
U5psfGRnDbtNU6o8hqd12RLPXAz9J0GJs8un4P4jZ3K2L5SEahW7xEnWGvSTSvRv
qAqWjOj/IrmAzi66hybknVsmlvcvnkiahMQOjLXJZKMQEeEiT6F4qymimY2iJLlx
GQ2PHz+PH+k3c4C9akXX51r9cEE26LDbPBmDLm0mBTmq5TTSIS4GyUUUaIHY6YfB
gvkxd3T9HpEMbd0SI8i3TNSKidoDa89LADQ9JLTSjeO1Vt3c9YZi2imB8u7XQgY8
lk/pLCoOoNFeR7AObg3/bBHpqkTvH/pj+0P9gw8QgPZJHnRpjtwZsM1+SL+vtPgs
Q3MzdtmuKqFdm59Vso38jlbUHDhGVwMfDF8yiIdriqN0PEo3sNPI1RQT6vbjtZPP
gZWrGuGdXUDO5hvdQRT+zfXKoMo6lSAFTYzb75iLRi902J2zMlLe1PRVu9meCqf5
2Ecq5bTQa5qtGjfB+cCYctIY/57DG84HBIWIvHfSc+9uszy3q3G4ZuGJFRI/N389
KNmlVrc5etNblM/DDz1a1e2tRpPff5qh9KIZKCRIltYzYM3XE+YVx02mEHTUqrYW
mfZDscztsH//+O+1XLGW8S0YqeXSXxS97da9+Q08MTmawvY2goIjA23IxJ9uC4GA
94r3oAGpdo7f1IVi7herlziQ6UMhzVfGOu1Vm/+6h507/FcV+2eCbLivKcJAibu9
X6S1RENvJ0wuyq+M8hh0Tly9RJtaXJTQzuGTbf7Zl6uUnYT/UUH6b8cPWKyrWpMp
nsJTeopmWmXnvkWiaKEOQ588CVTfdKFUuJFpZe6NG/HRauk4cwCxEg3yFLfCHZHr
khFjePOstzBfHuOahNoakEfutM39WVoG5NO8saKrNEg3i2tt843ZNKzf4LE9Rwf2
Ddem4Hk9ePqHXdfkGIzMTfWkVDmH2GmyuVLDIApNY7+PvilhD+0utR4xIf4GBnep
3D9QtTERzO+/07MWyPCTuj8fX0LzLMRl5nTfGkuIX69wVAjB3bEJ+6KfmDPjzfvw
lrZNJqzWdGLiNrVcxLwOnBeADq4Uq+jWH2ngGvDl6EF17pCvnQN6y+l0jPn23AEu
R5mZ7kWxsbCt1mPG/PkU9AE+qQd4aGwVu4yLWIr/hbWkb4h8y7xq6TAa9jChDeTf
WGcDsxsyseHXJRt+CrqjCxSVR7EctkNsRTW5lGj5BrylQ3yd/xv88I32cqVEVzLf
g2Ee4b29shND3kLueFUw5aJsr/1l5uqzQkHv+PTb+hncr4tc6LMAGuM0E0+tybs9
fQRNXO+bVrJz9TfA/BHxJEfQRMmSd4tUcDKTP4IZ9nPbSNVhuXZtM29tBAbriNmK
cgYaeZjfEmAepy1FOryh7b8Z42nlWt409V8n2chfZA+YYgkkJg/teb5Q09rFGVEt
hljVp/OoIrEiPKYcDdUkGwg64xH2MxgueGf79m81BNsdUB/LAIFeLudiG9dTDxfB
y4+CqyNODMLhcBRtKYk8SUi3AYhK447BKy9vDGeX4xh7T9Bjy1IMSzWHPwdlbCwO
tpmNcMVALw1tzRl4fuLGu2FoEqpSk8FJqMOew/DwynzutJve7OHPZ4AhP89es89M
xpg/85KUJWKEAcECAN7z2GwtWXb+Wao/2DVKKdvA1VcEyhvd+9V59vR6MUUhLwT3
50zulYs967lzCyNeFGljSMwwKYxaIvdQeHXWzMi56kG8bJR53djvg44mzgJcdYha
Bl6RLfcLQpENIVHcXeMUVHMaJmpxv+cIMhygvF7jLO7UNWdkEuRUIS06fRbmwICV
PqRXi/aC0t8x/hj+bNtN2N0kTBtpHmiLuCqfQdJpoVK+ljuFpBjUhndKEDNNZude
d+sFEiN/wHz2UOeDFxCJKr9oLet8AEAe392tIueJ/PZtPydgmXM1A5jLnr9OnGB/
bkIKMfTh2R9bGWffSNNaln/tvNwJJ2G1Lxdh0r3ocxmVGbybkIet0uqrxs1CXkZU
eFCHRIDT+1E1wa33kamEfzfd771IEjCxktwueBqpmY9DxbQN3jrRSzPdeByJEG4C
qMEsdcCm+v8QNC5crQSBAkf8HdXcL85E+xM0jgKQbrUOJ6vgktPAmHLbxBrTZwzJ
GWm6IX674mG9nkR1+4dMyBeShMUQiJFtIfmb2fQ9OR9vyP9n8hh3Ov6IQvI4shyK
R+95VZ0XGIQQ4F5vEj0+9mR1PAAqFILZdgjJ6gxMGASTjmPay66ASkNAz76Uaivi
DzHW1wQoKx0Pe9swhv7iho9RFCgegHZjkNza7N7t83UqTpsy3UHDBp1la5IDFCKW
JkQZqGgegBv57yQIp/mOLmyJEwuu8uUErXFWSBkEXN7Z6ZYp0JqQh+uVeCDvhbJa
zZ6ef1ZyYKKRpBB2srkkoPycLDkgzYEpbo9Wz5WQlphmXtTGlrzM6bONk7nftrbH
JaOG10X9xIedpG+Jn21ruIqtMYiJK34avhqpe1TvPFa85RTVmZFWWSmxy84kxfaV
fV7aFXDYrfb+jSV7v1yVs2H6ULCGrsRicCVVBgyPvD6UQq50iimKAcYAupYvSC5W
Y7cSChlLubGx4lxskV6o8jMb4/cpvQk1Ijq8NZRY16sHtUJBdY+bK05mBA5lHRsO
Q46xO6HFAVphyeBcC3Nxt8iZH2H1NL5kHxywLKWvyMTaw2duKcY349MGG8JUffiP
wqV+EHJyMX7npD8WV1JD5kUb6zn2QeBlbSEQDMaSVlU6s7vfSBmvM0bnOd7W0uXc
K+NaTDT1OpgpVRVaeF4wTt1KeIuJfDdujVSEyR3ddC6wjzWle4gFEfTMYO1S+B0S
dq0xRURIW3DS53ll7B07Ih9Baq3pSpwSQDsRbK+xs8/oxh1e6NdadgnjUiN2drxE
wT5EoHgc3gZMvygC2Ox//qlRyAHPwtmsz1LLSQ7xwMLQAQIJM7XHSrthvvTtYWeP
v++BIN3rjSGF3/mbrmRMHzMm4Tyy/Ev1IltVvE/6N4BJXGOgRKeAgOHOGbgCyUY6
fpT1LJCTbK0n4IHCp90NQmoBGq38SlnZQYxHShEXs87O5K7n0n6v6h67HQUz2/q+
B5XzJWKdBNU0eCSxMliGr7EkL8SDGT9P6XKvrrzoS8w/9v+d3qpo/9NOX/cX9Nxg
Z5ISJ/lAiJMqEvldG+lyRdF82p3id3S2TgSju5pzyFs646ITv89ubtItE2YH7PRZ
NfIU8uPNQ8jk5+ZOc1zC7YfEMRAzSwEIsdfCpfcuhXpD+/fKgbMONPwBwB/s9D/y
aVdHJvI2v32WN0CvxpUv0BQkaTno+hTAjqoP4+yH91iSQAuC+c3As3jO0gBa6YV6
Znsj+YPFcKHzmMEPqHei8SkJb9K1gIbaL+ZPFqg5UWO3GLUV/FrJTvTLa00LI5NY
GYWcxUbe4OsK+nxvURoDA0bj4EPGAAEWeoU8bPdJ5OLTurFFJwgRGSfNIhYGkqTI
jVD6hQ4R2q+JWqxswzQax1x21ceGu4O/fXU72cgMDwk9iG71851vZJ2eCz+nyp3v
LxMy2ylFTVtD5vDy0DxuijGE5RhDjGHOBJjLlQW5i2QysX8qB92bj4x07123nbbV
BFHidI+BvbNldu8rZt1FMXyfyzNkQl+ehJtrQrxF6ljVHfXJ0p2hecMO4gNFtFaO
mE2U5N2lIWWNDgKdPWPqzW7JsCWo67VkLgF2qz2X7GQU2JE9eIVscvyBEPnNt7Lp
KxkTmbVQndvybrQ6ZOe71V/+1pGdVZ1olBblu58b0bIY9AxYbWMdRwtFKl7P4vxN
Rqf4yRAJo+H3SN7BW/kUXcDs6xhhTXTG/Ql5GlilwR5rKrLUlgiKep6zhWwudNtB
YyyMC5XfMgN4oKrES1OE+2w2Fct3JuPjueXksls5NW5sewy2RGqekbgtaAF/YUgP
2iW2fG+3tIyJlYEpFgQLg5VGvELCjJiQOrHivcUnMPgbcwvTZZzx9EViQbxO+Vj+
zQgg9dbUcy/6ltDvDsducWrcp7bStYLeXadnektW2jaJOXwYphTO7Jasyu6LdRk9
ePyZmA0wjPr2BZNk2VAmx7RGRGKfc6yoLtE2QxXJFsakllJTdE7heByL2MkjSvbe
aLXqjPVZ6yMsoK8GcIRz2x517Q2pu0tlchESjXrICWYs7DJHYNVZsHEyHBg9CSlm
xgbqkTJo8jWjiW+UmkZc+y6w1GepgUV8LFei8pdCR6rG4r5PNGr3PtpyL0xfMIJs
6srcnB8iNWdtmrdb6njCz5ErmNiE5aMqkvhogBJvj7Q4r9sFT5lkX0EzBWzA6EEl
SVvAminlhXjF0jjGJPlae05XqPd5xvQr76dkiGv2t6OkbYt9UGsSddM+jgR3P8Ng
7NJvUY5mqTnlzrlmmrJbPTFhHBx9sOxXSQhPELWWsFsJMVgqkmOhqG21YFkTCQIP
yfmochJscp1TBJgFDRd9ZVhUzKW9asW57G+4QcJBvjF9881jPXr3/kngheuMSlE/
gkaFX41wBfUs4g/gAxRG7TPTjdp/zimyIRm2g9fCgSWSZ8nrW42jlHC0CFQ3mtj5
5AUI1umb6jr9pOvkEidYhydZ3bGY+sNUzM+JFswT66XUDa6xhJy7Q3E8BWMaDjjB
+AtoBNUDk+sVDq2XZGq3TjcPXKBVUEu+SHB/Vzt3iZnZ2vRE+R5BQdLsBxBhO2ZJ
1suYc5VJ3DG1Cr2336IMaXrepc62uUFz5pINuAlFG7plHg0wbCp7WH+kRRoO/R+/
1mQ7nQFCU2l8JRw6b/nz9zQ41HqHYd1oNXhZnJVi5YSpm51ISnllUZ6xD+O5H907
UyqzI99F4sghF7Tz2rm8g5so2XgCQnTDPkc8Eus5AB4uHagrhFIhVHcOOqdTs7vW
DFh4jtYbeWK/RNH+5ebmpc9hfwomgDj3ghIk8vdtK62pLSyKv5ztHaIZ0abbawpq
kVV5PCvgyCliAKpxdTCIyZrDBizDo/OGzfCLF3GCEsQ41kyz8mZSeQ5EYSdEJuNQ
jMe8H2owK29YpNvm5SISB/0OCXxjOyKmTXUAvTFjctfoDtRC+M9Ylu9pk0xsShlB
+Sc11M26gC8F5pQWixkpxnFvjt5aRc2XRpz4npTuLcaC+uH1mldD5NkwXID/Z5Ta
4O9OsBh6utdQLOg92UtkeLFd8FElz3vufBTGgBMANcvFlLi/ZioBFGvGLJTEWHY4
MFLU1ho2y95KNX9HUwWO7/3b0psqfosTF9jgAOhxmRjGkxf80Us1rU/kbSfuK7lr
mvxU6s84zLlKUAS06nzNm0yvBT16LsgHQaoONQ8g4aTKmUQ4O1PC2BEIlA9Yq84f
onQhMqI/FUubiAM9gr3bu+t0OLOH/yqyS0dbTqRxUJls4/2HAudw7lbS240SyRDL
XJOVoLRMW6n0J7bw3646mnQPzUiF1fdbAmxD0TWIngJwOuQ9HTyzsMXci2yjpI27
SoViHnmYieJ1qZOh9+/kl9uLcquh9uNxrmU0tcQ0THl96TAAe/EQERvbM+QpL1yD
x2YZEn7dpNa18YOqcsJfnKnrAbl4lNuoP5bLw2yqpFrxvpUDTa6Wtr999SQm2s3a
/vevqfIOir7Stf+R8pNG5YcxITGjK76zHejUAHWkR9/X0/diESFVaxJm3S18IXoN
aTUV8e2TwYUqJ6dCV2e4Ebs9WrMidD9Ufoy0fvNga3EaVGT+Z9HEPh4cw5mZ+OiF
mk2hg5Vr0PR4hpAvwQR/1L3XzDP/GjE7mwx0Z+AKLrTScQcWb+zLDPydixi5MYdw
ZkGJh5unQvPvmwgwH4CEfnMW7zr3oIR2X+sxJmGXFPziHRto4MxS/QS/4lscEOx7
+jYuM11ZIY39REOGfT+lpemIN0Pxt4Ml7rjCkfqATLp52sUvjyFPSdFtnHEj7O7U
Km23RE8da3xp3HNSUWsBF9pritB5o+Hq3SBmZn/55hQ4DD2bo/4w9wTIgo1DyUuS
EmJnKFctCloFH63icYK72aDuo3LFa++9pSrfuUPEo9rjvVCHLAokGoAlKujQKk1B
cESWsE8bwZu5InM8FaRFBMgF/Tb/Uc//NnhdgCWiwB7AfDHku8e34MX07IpaThhr
0iq4lZdMKCDfq7jnVHsy5RIf9fPmHPzLKe+ZdJEaprq1CNJTIv6QekphGjYfzQM2
TReYWc8aNd2fP3hoy2cPa/KJFiC7L4AGb9mfrRhVRXj+AmNuuWuuEV8N6nam3iH4
LyoHwSkuk7v1FfSVCBLn/e32KwSbcXW3jzDKDL/hyTpePNvMH579zaUWzHNzlnsP
vOv116FDI+T23lkd9OtascTqAIzC6ilImTlviN+OSovCzFdSTJVyfaLYD3LxWHuJ
Y35XuYvhXX3p+4otnFPd3iURzldHs3IJ6g8TSMu0U3JuWeqGS+EFpjfAqRAa9dbz
01F2GeTlUNDU72lMk9K4gw6XGXsOQ7EhwnjaXdAzdyOLbPwqwsoqupteuMM6IsAN
5XUblWoPrFqDwl/2UYHcRwLva6d5yyfODI77iNT9lA6XZih0HsM6Rl6in5GTUiis
vie+DdDjxLrKMb22X6FAkKh2yyw1KtdXLb7eOI9n5KnUG1FkL4NIgA7t8VI8LlTk
nPQpKdP6t4Sn1vN10ZDsL9B2elxt9eZVbxgYwSLHp5+QdkI6EPWnvIozFflTUJTs
hq1vx6AV3BjfCN/8RiOYpSkLu9XlawhU+n1Le690uKN3X/z0r/xAev8j2CpcyRYC
dwd6J7OaTNyYmzfbJuwqMW9ZrH+miYb0FpCUPP74HmWplCtsNqBA4v3qguFyGtP8
TxoTfFqeJusSm7NCdSKoHPZiddfZR9FChV9wa1wSixY27xrsqgTVcFe2G3MfMi0a
WcxeP2c8SVS7Yq09Dqjw3Wh8ZZF+Xeh8AEAdpWXbn6pZaDaDe4PxHXBhi8gd086U
7PI0vFO8H2ur7A/g7vPyAL1RuNWhdld3va3gWmyBU/lephK8fEZ6qmSZe3Htfb5r
EsZBGPPJfBjCTeMRyfZqLcqMty2Xqn7ICzcMet/8I2UTWjZFVYFjOwNV6/GrQHKn
wqTnNzMxp8u7fbccxqdPvks4+d2eu34MEG3Zob/tO4iEYMdaLOhF6mgr0RkdQZxB
0HGVzRl+RmNYDvdRlXVkJJ+4RJnj42au5kDH41lZ+hiBFVbNxDh3PI0XDw1sbnbh
Kb4uf8wKRLYqLDuwFia68awBI+9TuhCdnkyQN0DqOohxtlQC3cxrOHd5JPSm1eUq
/lEc1H7i0+sgYrdMrOInS7Fx6IyxY6RRELFWsL7vErdjKio7mVijTuIiPyUsFBEa
qlMWEzZk0nHKyv/6DeCTjiuNcCv3PzYUuS8/4R6kjM+68PhbUgI2lwV2Z4+slkru
QrkVYafNn2HSBQReoNExsnPspNr6H6wZf72GKTZaFFUWCOHRd9WR/Ky+gLvbK7Sh
IAAGOHXiFDE/v7/9KE2WD1/mFXPrEw2bSeLjcH7Afi9r9iBHNpF0+CD9ONFMupkl
6CLWIWb6TieWeZ/UYkQnTjuXhH8Uu1lJyKsrVb/kBiIgNp5QOn5VTqr9yeQD0LYu
sLX2XFp5t2nlt4uymX7Jfe/wWK6wsFS0XmgJ3s4lmPMXNiKS9YtEQTfVRW3HoOFh
eSRGHIt61dyDz+ZE2goz7olqeucw1l5yjMcrUIOuIYe3PseYnEJSAPgb6dWhheOG
egsSXqIqfH+xDX8VxOhNwNfWGHHL/TUZdl85fuEs2ZTD4AdQjzKWR0pDMIoUZgcm
gCDnSqBMikEoNjG5PaF5a10KEP64Mw8dABISU9WYJt/yR/+0PnyQEShdlDHjohLD
smp7X2n5g1i0xmLDvtWmpFHf5LFgUaSzAUX0Y0eUE94UCqiig2GC3xhAzKE52fbE
h2rXgl0WakFPukObnQ92RO9I0Q6W3rdnOdOrDXfD4ELdHvdeKGrQoh5bgrCcAT0o
YMFypO1LbWOJMWHrFK0wlzcrXjkAmQiCLFJgbGwG5DmD8sL2bLvEcmWOPy+iPNxi
rjEFR/nbDnr4tgyXQL6kO9tiQAqiaDFeK6pSRgAjqkhfjGX3SgeK1rebOBv4e2Gq
LU8NiT43z8iwyTNJ+QfQ4Vc7DZhEq2JcQWp9Q5vch5y5KY3q/LJD6LTRgWkSnFMn
XKbt36YB3Lwu0q6ut0PXmGF2EQDp35dh5b7my5piS/8iLI11Fdn0+tdmV1bvsesF
kCThn4QBL2GGuA4+3Tn0mIjOUREhXPjU/BNmf0CEpSWWJyqQP+clpcy8lT0i2oKN
EzUQ52WJfr+HSLthPGtphZ2TD9f5QTObCD7kQ3PFxhfkI582znVigVRwp4tfAbbH
5Jyz1DXyMX4bmP+fFcjWVsmgaS804j686vCLbjJ6b1WhN03Bl3PBMMykj9um5vJD
oDf/iLFPDhMVlErfVGUe/8xGebZcwSvpXT/tm3/rFhw8PH1WF/oy+qXc+aFUIEGu
6LAfvmVbpnw1/g5KQ1g9QfSxSAcqenaULOShgWMPz2f4em125WS/AAWHStkE+YrQ
vznB5OTAXjJlPWtdnpoguU2Gz3DeU0zwY9f4tqSFfBWXmQPqwPZavFdYAalnP2oY
yYf3jsh9ASRYy3nvGKbmObP/d+iiR9AQU/IgbjSDVNxEcjiYH9BaLWMv/nkyIGh4
GiTWjPJbId2YS3ishmxPHOhejkBwfuKXI4lgMryKBBLX0xUarixYPBXm+uHBarT/
1glo/oPUqEBP3dqSkOK4qp7Ct9j6eJtMKn0Sa4ER4vGTO88nsVkEM3g+Zqp2L2lY
B+n55scoH484in6DyrSnxI9g+ABb333RalciUyDVYJM8Y3Q+A7Wp3clvDD/0m8rD
xzpPmaYSaCdN/BYaIWoa3b7h6CEis0cyVhXIITWoPFFU3yO1IEKEZdIgkeg4PWBN
j5EyNyhfsfNbBi5zDBFfVGUn5lhV+VLunYENBfFAFobTByj6asokIoh0JUKwtk0G
KrZmNgHyNq7kJB52Z7oQdzaJgZHNfd47yplj3Ysz10gBfkKDjoh+SokuPAJPFyUk
uhpzOilfIYsUoaKe4zcIFFLnAG22DcydijIW+z/CkQIULf9JTMsG69E77QDxAS8m
xpaIAGxJff5ABm+boK9cDCLBnQv0BLaZCsBU7Fgpol+bcCPadpOPOIy2hL73jjvP
QOfQ39z3aawfa+AWl3C9JtoSb32UhRwZki4xbWrDPuWuXwqyaDjFLodIqwRm6YmB
i356Zfhqh89jNgYQVyPypsKw1YjoHM4WTP5GbMSyI+ID2DbMKIk4HFDu/aQLfprO
nRxG8Cnkbx6/PCXFiOvWfMXOcIr6MhTxJOF+MR3iTms9/DbwTZjw/rGOaUhe5t/Z
Z6qUGKN8UTeM7O2/3kxvJg934xRZxvA+QgzhD+X5WUtDM08phSwMxAPa6JeqTO9S
cHLNiMSGW/l6k8PGiVrYv4ffgRy6VhDOBB8ykDLW7/actCAsni4Nh0nn4LolB8rt
dxa3m8fa4nwFBsP3vMgI3k3oLnxDghhFxYl8RPUtnseG3/7Zo4Z11NHYnlrk7DMx
jsuLVrBhhEITNWdq6dch1qAn0wRiWlTI/0+u1LzWSfvu1PGpzaLRm3lVVKdaA1uV
0qYT7uolBOdQ6Acm8ucKFwQ30jhgxm8jAbxV/9jn8wzfGpB2iG8leoBvYBaVQCg4
gRoZrbm2wbkwlXqpinymCpPO2yHub0xffa+5lYYGm9MlDxXyzTXubANt8psRl4de
r3d2r1OxUt/Uhxc8iJmT4xXg+Vpt19M+lLz1iU98uqld9WAkbWL1A5hNruOlq1yb
+bIgMU5WymH65/1qDCj6W+DajEKOFCt1Yx2D22ZAjpthbvJt0WHoSlwud8yEwZIt
7ez9S4TsvILeKJxxAvBf0v7qMcp1hi/CxAJW6ZJVZOMykWnFQcHZo8+WkM9uPNRj
A7IVobnsP88l74/2pbVRW2iJhWEOUoYtuye2GEZUAbzw3wv2xVZGEXjUZqNibEJX
gY5UgpKjt07xomkfwksE091lx5AGyUwbgaiNSvwEKBHlS4x89X/GEr3L4dvvOiEx
Z8TqVeJAx2GJDEyFJ5wfNOHWEqc1dlYowZRUYDW35sMfZ+dxMMupMOc6Ty71+kfR
uzHIsPoBpxhB52r2WLGOfp6hbx/NnEEycBfGS8T2H69XILzJrK2zPu0tIwrMEa0e
ITzwJ0npGtJqlXI7V+leyxW7gqP7DIcRUFOeBKTtfAnZ1SDFcokbe4vrzp1Z+4Wv
IHTA11usICIriyVfOkHrBKLIUaBVZRX8Tgmfj2/4/O+qPfzho61c8QBVvLXI6QKE
2TiasDi1tc3ZNvo8kos08sn36k7ohOydnDm+RUcMMBgjrs2a/wHQVZjch5RHAcyB
NlrV6zqCleLcNv8o1SRYd42dCI79OsWfL707MHojbAccgnnUvY9ia/STAtuza2PH
jg5HVUoUy6hv0B0a4WsEZWIPKBG8yMH9b3yPkQKknN5Jx0YLfN2L5BGun3/nd0fP
pS09N4MWGTXcNVOLooj3z4sL5KoJl3M17nsiQv45jJUapiRdhrzg8xxT8QHMNNj6
Ab4OXsuOeGKk0qQBoYkgwgJKIkILQTqapq07F6xa9oU2KTi9V4zDxsdgY7c4vN4X
VjCO+s0rXgSBPPaUVa4HtkTCVRvqBfV2BzO8psT5BlYWMfyspk3z2rvrpJch1oUe
rGsu0rbuqyIwGg6NIw/PixWRRmTepUTOBt4/0LUHfP8LcJT63JXjxKB6kqX62eNG
run/cpgIm8vDomSp3uJuQRCvYY3Hep4PINYJ/28lM2+ziEYKw6WWpgd5lRXpr5t/
TI4maZXl7dzfeqTjd/ZDpKxZAA+KpbT4qHp0LgkyPslCW85C/DhRBQZQ4fyx+tra
HafyPECsNQc50q1HaPOeruyT6hMJyoMQFCUa4B+seN3E7421lz9brTFMW3ZaVmSw
Yg9iRdqN1LFlmqQ/vkYq1tv6J5A09iPB2A4qTNZ443PfGkgXav1MX+QLEeNCS3hV
ir1iQjjIFl4opzvL5qQyepEH59bgk1A2WUPOCqkjGl4H80MqdokcAYYuecKdF5Fw
xgyp/XupXhNyvPjNOA38SVYYyhNOClOYXBgvxpxJ3+GceXo7Me2r63rkEMBTFrV9
p3kkvm42PCnCzHMxkQJPCZtS/FXSFuC2Muv94+NbuXk6H3e2KilQMNL1Z8mbExix
xkkQvZ+m/C7m357OhN4Gw/WpoPeJ7VZfw0F0ViV9o2NMN2aiAspCcevcK6PFEnt6
aSs9qsavdClx1rS4VwJ/M9za5oR3r6AdQwTAJiMv/k6EQc1U/xnkL78OqaRQVAg5
imdgHi+6xMZa9ddvfetglO3qmiCFQh+M/kvMrZtZ7tV1gxGPZWQZxSCOaZKUg/Ty
hMkOC5UcgYAFIoZWVjkYe7ZcdCSbhC2XcmdTtlE6rG8Aas1+EsGFI8qnA2/HF0e3
ZaoeQLmnDe/9yIqUMTqfMRfDec7kUQ8q+tbnMAA2NmOqKh181lmUCIiLiEOrYiqe
4eVxjMhekflWBp2TqpJi+mqfloM7mSdJqh4AjQiNl9G0W9f4AKYMDD142B1MUxFk
bFl1pMeDypj14aRH5Oaii5QUbo4ftvypggoy2kPywmHepDuWuNHw48l/gbfbqFG+
C1DrQ5zpIKk49Wn2TPcVyvs9K2kjibEFRrFJp08zbQtr7SGWWSHNMuhG4qFJCuQM
BR4T2isxBBWHvlJwdxEXAgmEg40MotLRM0qka+oh2o+7HZ24JuOr1/31aM3o7our
h1Io7NN3h22GuhRd7Q035tDW79dNH8vi7MpPZEZ7fFHih7wDZfPvMnqDFXuL+Hdx
cWhs09xgKuBkdJJ9dzOGqfgNaSoBr4MXmeADZNFSAsr4/UnJMlFdquMFjydxsBzP
+xcz+AE7ubWnyyuQOVPHOE4lKRbl1GKKgYIiePYeR1dIPAtiRT4chSiCMusKHDur
4gVpohbNUKAluthPr2f1aFbEtEvQguKVT/Wjwmm1VIvnkso5ziLl2Ze60HD6NH4P
tSuMYqF58YC/JL284Cjcf0cZBe8XVYas9HYnkY0BLofVY/7uxKDpTqP3ozuhYWhX
a1GBrFrQYutvvF1iXTyqdrH7eDxp+EdO1Jn74BZpB4Tqlx5I9cP5RjeJm01pobiM
KdZEY1LZApLk7hKeabED6fvgmKX06DUQMQllATKvTs4P94jXdzLDRyreLmIAIqOR
vbruVJMccxLqN9//NBWyF8hg6MIZqWM9MtrgkFRpQjyK2REJ3FPPAH1xkkG4oO05
ypKHEXdQTxrbAj1bpPFZLG/QcbrpLruxLnOSMI7sz/6qoWVNLt5z0j7lLSyaRQ1m
nJ1o9xsCPUQKgItiXi2nvdSzr7xaZO50amBdTGvmlmLY1lANJ4c/oxeT1kTLLZnc
MP0Nm/OiJJm5uNVRq7F5qHgXvkMhAo4zYu0yv57U14qNmzMrRuk2hSscAhfEFu24
5WjpEULWwBiDjCqwDrpHuRZYxCwoPyX/yL8a+tGAwNmXkXERGE4LjpB2XedD0ZS8
e6ECgCo96T8MCH9r2L7ussAOv0Snw3I5HIZ3e/nx+fnBhV29FFA3YhvcCg8Uoh6x
r3ZknkacbJ+eYRiiX7RrIW/FUjf8p2uAHM9+ST3/nMLI1thKfuEwU9LdzX6LPCP9
jjzmAh59Y8O42h/r4MdONksZV02MCRtpnwayjdo1h+G/jMzTnJi6PWsURcbLtPWM
4zH5VPIUVC/IG5aPC8blDflFsGjDL3BOY4U/NNDc+ZONf4HFb+x/y4aCLwMiOqab
ILXZVrYwuNxHxOIu0K5qLzN0e/0uTwFVYBccZ4yhccHlXEo8AD5J1JCpXqPQJfv7
b//ur9vK2M1Any3sP3Y+z35S9sIdsQ8gDtVRSopuTzq4Z3sKbf7FqO0e19Gij33S
AuRheBTkn9iaLCd8g4iWbnVFJxMAf3E9ozWIi+4biDVYX0gF/0KKD3TLK6RGPR+U
d06hu6aFctsQYptjQqG5koURa2Akoyf8t3euvV04KMvGxZy/rz7pwb6zMCz4R08/
coPMmD6MCpiBixr29LxZNXHwnx3Wg84po+CGNYW3anv0pNBCjnAM04gsmDcCPTYp
HG18SWkp8S4HXCCBvBXQLUVbugojdb5aA1bjRr4FD0Ezq58j5uBZb6BEyWOowPfK
oarkGyDNVSjrJ5wxByOZYgUW/6mcmWiVSUmAGqs9EpbVVBWe0Amej5T44VAdOI4x
pXu8HvXVleUwQ8vY0xbANXE7ca02Ia10ZyPld09scujQLEzPuLkFurif1r9dC6Zl
L1v6yHACmi/z96ZmQenbkvwSml7HDTiadiXx4oGGuFBRzZu33cNt7aRpArFmQ/Iy
aGJRwZhgLl6gp6hesiCVSpJ39NVYNU7HE0ut/s8b//IB3nLoQ/ZouRgZd1OU181v
m/mwAOP3dV3dPjZ6hCmbcygoah5mwCzVITvz2W1zlZRxhp2OuSzZSVYpZ8LKVq1N
5/QjARu5cETmWE8HV3QohorRC2iB6eVHLDx6HhKLjCHl2B/w2FJzFC40Mnp3lSoF
ceCg2MzJUZgObU2l4V1QAxIz5ZPV4V4Am3xZ7Ct2tnSMvtWR+PhRSPnoQlOBSnnm
RJBeix7ZC70dwbhrpp9+rat/xzLqsjcmLQtsmhtGK30s102VcE6MCqci/blHF6pY
/YBkBHxRIOOEZ/5oZCvFObvNTYuoiD+217Vs//8vsswWqiDT9Jh7eXDPRJrm9G4G
3uBw8tCfnIo/DSegQMC8PqZ6Ax72JB9DxSjljawd4yWeGIGGwlMp709CtVFzhgLG
pUWZ/lmJz7FEzYyqC9LyJIbtzVlsKXPWUohKOzBdTL0H4rI49ZES0PLf0pKNh3Hq
SQ6sdpe5fsnDVb5OMMLL7BZU+qgr+qzQ/lj9FTBLxu0ITXI4jFXpM4YxWGtuFvm1
I7om5T2e/U1GElNgwVa4xvwponflP8Ln7BXM0vLFdZNTR+zXFL3qSb5pzKt18M1u
BQOzcBaA7q6YebJduZx/imGwXABdOrbErxf54gmjja1BTRMSYrHj1g1pWNTU2aHl
OjinQVtFHYS+Y3n7WiK/s894z7+mhXZVJVY3q2jz97XVTs/XrRXyjBvwTWA5t/Cj
Q+lZ0uWAq1QvFWMNrqyD2YEFyGgu+Osa+MNBvRkrgvYnNqj8JGouapO1DEpUhXt8
9VCvZYc900aMF2embMUE7z9bnioL8iWcdc9ea/D0hJZyY+CjVsxwbAehpNgidSGI
GIeNo5UdTIUq39QOPjEt5QN3dWImb0TFAqLgjKxiTxwmjof3Kknkgk7fvRekDHF6
o9exSU9AC7gi46L0AH+TPxnWL/c6mP2Ee99G2qrUZeGJImdJ66ePwuO2vl+Ei4Rz
utLdPqN3wRnGi1uNLHY8irAsIl2vSBbjUN/2GpgUE8qunLLldTHKwpKcioIApNnF
GbWKvPK5xiospFQUdDM06ZURK3dD4U/WIMDH3u0Uwfs6lT+Nbwf0TbkIoiIy8tEP
61rgwAFhibJklBL1mN1W9fgtesLSwH72X7k9uqcjqHNO+hgE9GAZmdyZZQbWmUzT
3FwNOObuITERaY5Fv3ONsRE95Ufd7S1VDUaCA2tBQb3/meU7QznFks/0wuxOYtZx
akqiLlMIOjlbWaYtbN8BFsv19eFeH/NmxCU4f+ltSdhqLfbcUypcWnMj2T5ESjmI
S8WHwWSn6OoSU4cfLRSceXX1ztuI4fe5Yj0ZV1Ao3uk/c14W41dNg4fbKp6/y9KM
1J4sC7fNhuygpiuor+bYn2JnMvDJ+R1vz5jB4wSeb+IAOOwoPuMzj+zcj5hunxPc
eHHH67T2kgY4NdeXNuWko7Y49JdZrwajLoEkCXqlWolp4ZmBwKzyWBb34qS0MkfG
BelEzKC119G3QzLSdP2h8xLeQ4JMvHwSIHgWiUETbYVPPQ6+FejNHwa8vI3N0JEh
1A4jg9Z36QyaeWdJMMtqDblMUX1yYjJZ42kOAaKA3B0bUe2fec7PCssXBk4NAg0R
UhKkNut1LsteM0nAuNL/5LlgI3A6RYfHyU+iA5uXDg7Q4Qupsn6lyJRJgiytK3cC
O/fAsBd/hIJG7OUigdyWIqqBIVpm0AB29dZB3xW7wXuEdsD54cXcC0DTVOFQ46fH
wubw0LpnNH46yzr7V6+9wL8UEBTZruLqZoAfRCDoIiH3Kj00tjGJb7JngLN6IfpT
IJ2H53E1aBN20aoTTO3gMyXWo5Qjn870OFfgYNa0ZIpwloTU0DYTjBi9bEiByQfW
hUhRJI2ushs4AK19nGEUEkvul26aXVTiY8VingNMh0xambWwRcmQKfz19pH12WIn
e/8HI2/oZhnfYs8i+I6njqjz22QsaJl6cA3MTbh2wCdVNKndDwbKVG35XswtnxHY
ZSY85VDHwZMshLkOj2XMPSxnHZNgcCv86DGq71ZJSGcxwMwWd6d5pnV241BUI70S
zPB8rdXCxWDsKrIjfB5tb11pC97Z5AcMFoQ7le41CJ9FXTDq8XKH76xpjozJRkJX
rh3EvQpSP8AKAS9FYlDLjV35d7fQsU8q+GhDZ6TAsrXWQZVLpfqEcIJ04fqwxw6L
1Q6kCVnLi262DFu7hbGmv/7d9H1SVyFPTItecSqEFgTkpUXQJ7iuzdAJ3hv15bRG
zaj0MhdM6pquhuDqykMTqO79zAsCHQwjnNBR4+AdZHI0ykMJZ2eyYN+Dt4LZbKUK
JbJksU42Zn4LBogD3mI2dcBDAkt6PecVlXjfOkiyRm8dSohrEdWPXPg7OEF7p709
tOzeXqPQa/l+jjNhikmTz1JibW9QoxGq0EaJ0nJPESwQk3HddFk5f8+WXH3M2jty
Rnj5hSM6jqHMU6dsvVPWbAIq0Vb5fh0VlZ7mUr8WNfJpB2xhO/CWhg3LzvNjaIzh
Y4+4kLa+dwS+1XDANoeQMFiEJGcYP6Jy5BBqah17BsrjUf6XgyBS8KBfcsJaQMs3
Vp7NjfkVBAAxl/I0Mn1FPYIgrf0RtFbr8XEF6E9u2BHb2Hb9MdhX5Fwd3zF9MkvB
WU3ASHqU9vtyozSRDCsai2Xs91HSOD9hTfb39P/Pv+FFmEPru5QqVHd9vvCMS3+H
WAhiqNazYQL/YUGgVYtOxHN31NvrdKSjwV+JOgiFpwW0XCLvOV/JeMoe5xyTDBcx
NBW8EEM4lyoA3gMhvV85Q7uzAFlf00ZMUa6lmrdgPkMDpLCGYqw2P61hEVGcRJ5x
oM3kvGVxh8F7Jb+ZYmmAwrkVIJVRbOQlx+aqhE2/Loko8myMRHmfEJxE8eQTbDLP
PbYmSoPs7r2mQ4MQ/aaIY8j5Tk8pGeVcIrTh7CD7nl1We4PsVCqwLv6Wv+d6FFnY
FAWn4BMhFwoCABynkkjAi5wuxl55i5tCzC/44HdYYT5mSRt0queSnxu/A9Fw2a3Q
acoz3I7BlXVMzXUoMCnLvBuZOnp6g/7C1plqWbMO9rFFd3MWpOpdm4fzT7VK/gMN
yWcXt1CGk62631xTwXVT5ByFl8bXTmD9jYkldwU+0QwVrreK8+smTwO5wIRH3Br/
2Li8pNnNLF9p5DyeILjmihwEwymFo2Y0cErX3SrFwlsCB6BE7bSHw/Hhg+a1QTaV
OrtKlxTqtjvoyXgR0+LAjrIy1yU7N932DMJQuXZCaXLloav7DF99kiH4NCmTSoo9
I+1+e2kSVihRDKtR/JpP7kmox6P2QzlYLrMjvRQ8AInlHSGIYupkVC2/mqAxDmP4
qG5lOfob/JVElT9JkHdF9D3fhJ7ldhIMIzwElMtQ1nCVwhy70m1FsRf8D016C7OI
Eu1ScEOoMgQ2gu+ldrWR783sZ+7SI5NWvg5fI9tw+UgfIe5NW4t8X+exry/q4EnN
cL/VzKCFb9GW5ZwaaXbSovEClljTvZFweqwWMgFKtL8oihED2aQJ9tp4QEAACINs
zWwNtzDDTFOapwRRrBURnLOa5yzyqj+POVqgLfssgP27fSbPNnlnH6V5Fj/VN9zv
eDhgqb28Ul0yDTAuq4DI9ImaOJCK8TcRmlOFoSRdlnCEaGuWWOKr9/puhAe7hrKr
L57QyyC6vlpYLLnVLQ8VqBh7yvwkJh5XoK9pXkcLs+a0NjIcxTDCaSaDdTIX9NaY
DR0RYzGd20yEYEP3y1k52KVHRPBm1dYD2UR/OzvL4ca2EtOwCzCF4Qp0dicxo9ni
3whFyn5S4kCTLsG1Op7zRD6pWe9TOtP1hJmORu8FV+c8BwnCGiycEF+bxmQOr15T
0pOOf/1m27C5qqFThvgvua7jPrjzFN2VVBTaLO883uGoK5PecO/3zYXVMXtMByFQ
lYvwc66GogBRJuKpX5g1PT20+d7kjBr29o4keGHgUNH4gcpTpwIU/ZyhN5BXnYgz
ZTvFVCNs1aWsHTQppX66l2d9C+MV7pbKvk933Qx+c2X4oxw1yRF9RJuVbzk7dge6
GvUBJ1o2SHTjXZj4PHthMwKbc4NbIz8Laa99Zvv+rrgrHnS77omqHYlLjioo2H7F
XpCcVNGokRcWasbHMor8bxozNafBLuEZveW+lq88Avb2jdGjGZIcL8N+cmPQK0NF
yEFyDL9Wqcq4oeKPjjKMORQ2azrFodEnlRGqfhIDjy9B1npuZ0PV3xRxSD1NoA+C
v/rx8lvTA6D8dhODcanQcKAOIaSwDeRXzK2GGIbN2BoZvuXXiQObkG1ApjZSfCfm
Gw5iFofy3eRkLbLg2m++AOwnrYw5fFIEHZf7Pg/fO+1G/3IvW39YT3/wz6myEVH/
vY6IRWVfXzDdqEmdAxeVwz7c8ZclLiychf2iJ4AOPD/MzreabHs8j7R5eBGumtcO
bEU6CbRl6RhbsIMFH/uocGNZ/KOVO8euNMLhdHpNmHAqFDIRejY7uBDPP/XoZ6Ux
tW3wUqZvaQKU6j1v7qJauwwfa8iOrtqX3Opw8fS6dR53EtQPh9NZohiie/nm2StN
9xgyeKIVe5H7XmzUGs13dxGf4SWobZh/ieiqDdCDGmiYhbkRJQCzMUFUHjUmSf6X
jn6VQorHYqjU0Sp9Oc+8bf+aOx9fDyl9+6RLTaM4lWHhQyKQ1OWDOulvT/Fu1ht4
iQfZx6sDOZdBKxbVI3eXgQ5FOuMhM3KZOQDVbpE6ka/k8oXog3x/5iYdvjQ3/Lcs
l1OBUWHKhvon8pWaicuvoTiwXz2qPivKG+UZDAMKR8pm7tie6Ew5cmJ+f1AIzyb9
BsnlASBRYv5HRq/cymgDNg3iuGrLlCOi566tCRqaxvo5JzD1jU6/2xx8OoMpmSOU
JNN12JfcgceL+FYSKe3oc0xZDE7ZIsB4eJeaaz2dsEve3/ElapVdCRXQs1ro4NSF
gjn+6ODZHT2GM5HhXLIiQ7F8K57wELqENC/bjRvLOXpuoYhn5UUGBmfOsf9HTPvK
xIdPyDcMsrdR1zuecSfFjB5yZQukUq8BN82l39ppygpkk+B6dVCurisq+v4ioWnZ
xMryceiYofR0IwXK/xsupFfKnyAxipaLdOct68mG+Vi2zfVo9cBhs0/5IDimTLMO
tmGOS6jhl9a7mYgYorLG+VGqbHv/t6zG1FGkHgDYeD4A+DKJ7IWQd5sIZywAdXV6
GnZZrddQhk5qzbHYIxUigSl11FY2MnfXAL6iunI7mS4AQQ+nPZ6KVf/CX/RxAOmg
CPBhC0HnQ2MKwqslSXKdn9V+JEMbH2hnbxj48nIIYfS5w/R/l4Iw+O50SU2ZHCHl
f0eFNB3t1tIombh1U5Mz0GG+6HX2C4ekm2ZxHTzXgapKq1yN36WUD36eIXIByAS+
Gam629yfqCdmHQkJE/XA2UWvz5Pty+dTfGaozsRWCEcEHbYpYXxAUenf7CvankAk
xjwVze/dJoPhRviadKVa60OIioTddb9v0hZu5l/lWxPluTEWmTe9MxnAOfVevVus
On1Ju8nJDDJBhipEJdrILUlpPFsJizuIeIJWRqNk78Z3stZvGPuVFO4iRxc0r+W1
sKSkbpJ5oz6J0zdPy8cyk4CRUmurO/BBvZwJuuGq+BEnLTr4mMd0PtNx//CI5cSp
4Br/kD5q6UjzvOtph45lk2bl0VPl6Aw9C3T7HHSV0fU4ZyW7Z2TqhJpmJwS/aruF
TFxJhKznsVf+Q2zd8tyon0e370jWEOIv3FEp/Pci3KiUjGGdudVuHwE/kmBUwBPO
/KvesKVHyRj4EYgmyNb+Yko3VAxMJT3dg4Dey9PTIre1a937w/VzrwV4Lj1aSMFV
VgJCVxKGhSlv3Pxnb12fpr6m2KO5uWCAKTAU3jokQqc/gt0vhsIk6GytO1+gIwlS
6j73KzZJmgIsr8GIpBB5Vax8rffRNdHi6PT7RlCsgsEPRAriI3i8Avvcsrg4sWeC
x17PIHU2UXgTslGza1xE6N5VorEvabHwY+ULyRZewrZl8Gvw/98KV9YfkAoHodVP
00588b+P55dO4z/O8X0koT02nUFHnj26KKSPVKGWduWFh0lgbSIyC7WR3lzp98rL
a9R3ZH2R4GK3dFn0u5d89zgtInZE9EumDTya2D+RNQULKA/gL79ySDZTR9EMsNEO
XSncsCAfycu7Yz/V41U/cDlzl3iwOETcDP3VIJyYIHDZl0uej36hzf0gqM/WZwbV
i+4AYcTV4TFtABcNaXUyQquraS7dFp+rPDt9izP+3iOm9LZFc2kN35JVVYtJd0vb
JtKDeYpS8Koh4yX6Pl/vfxlqPEtbfbvj9cvV39nUxA8h0eV1jXhw66h/xpt+XUFq
Av+mQnjDze86j9bSkJWJp6+CmO9Cca0Qjqm99SCNIz+DTTlGWbrtixiyB/qGEW8e
/JWTmJ6ljdsIEoVyoO9+gRsGPiMbnKyELu1eevmBTN1JNpKt9/n75x8awFsaIMEE
EvElHat65O5Wuo4JrwaKZqOKBz5FWoHPQd/HUWjwDkV07Z7auI6c8C2h4W+STOm5
FCDs/3/TmFyy/i2LsWj0YHRjshWbLzK5OhJjqRCpjjNHx68tEAwWejBQtcEVZEaF
uPVMPpJ3DsyZS/uR8rBwN+qt4Jos3cH8SzCczv2Z0jKTdcRtdqOUokqwPl46q6Ax
eDLkteIn9MZongnQoTCTWanzZ8JYDEeUbgOikq8eHlZvOWbl4MaYPGKIL5tZ9Zx4
BlmGSKM4F7/1qWxrU8LoSKeWHEmS9U9pTSdIRSST1Oniwq117yPtleXKRlHHkQgG
/nbLuye6AKG6eIt9btix1R/nUGz0O1YMB1rjhl/0QULxI83Wdj1ESjSpQH8Q8Zz+
oa6EixSpFtbyTNtU3QjeycidaLqWknx5lvbSDFVvdpdygaieDqv9YIbzyKQ9DGd3
HSgpxWZ1t9DFcr0wX+XIAgYRR7PVAZKW0Dk0g0UFWRWOjRnpl4dnzX4IJvSzCzR9
/QFjrTIgVEIjYj/+brPnIIBgFL8uVsvu7lWqnKB3RgF2ojiooMNUBxAOFf6cBjGP
iOBr8ROJ58UZ5F053XA+kUQbbzL8UO/ARoTopOw54RoiLZzLZ+iWFBFtBbye1aXZ
8rRTOra9ztWb/tz0u/ayuVjAUNBfXiXAbifqR3uASUkhoPYHRONYGf+YIxtH7TQI
h5DPn+tt8Fj3L+fuPHMF5lLPiTdH0+B+/c/UsFxJDLha67CC8LBVmxtIwR1QBvdH
37L8Ol8+bXycUuzlQE07aCDPVoHqrm4kXjwv9Wfcm1AIeSprKywDMuZFoJ9Xo63/
Sv3LB0n+YUlLAbQQsioVsOSJ5hZckF6i3oCSM17WvAn9LBk4MU7RadewksMQ7O7k
zTixvI8I51fSC4TrZbrPH2R2cQ7T1LBseTsJygdCJ8asl9sIJfU4zz/iwgQsc7sc
UV6CUUULYF36qy2grV/vbPkjPsbrd8vD3ILpc7VTICMuT9mZH3APokOOeCzugvgP
TWDzPwBF4Eg+S9wB6dXt1b6v4R1oL1D4UCnEitt91Q1iVsfYMfgPUjHAUwjYBAZt
rsNLCL8Ea0KOEkWihnlR3By7uTRUrs41wxegmmsE+I86maBFcOQnGR6xb9Me5yli
x1TbhxnteoILSEc38A4lr2FNi89H/9gBE1QuIysHGxy+ybXWwVAfZnKuZu6BBbbZ
+lYK+qAmuQv1N6bBWR+o7XeOpfT8vaTo8nECtfVZqo0F/6PUY5k6p/yHVjdvhLxO
WOVL+dRjHhD7kMkxcxWOyhLruubvQG46mH4n4GXKUa0wowPMz/x7HV0d8Q7808sy
zcRcWrzVKiXhWUOBukFYti31UC7jvRbrs6XHDgl9/pYNXffT0FrFJTo5OK5G67pZ
+KyIk+CVpcNfcifTB+YmCl6xxzxmZS2tt/9pX0l9FTp9JdJnnbamPG9uQaEUkfu8
WIlqiz8Mwtn9pVHXL1xFPWob4m5ZWvkNB9duqsmVUammkmomAEho7CQ/wQAlkP5/
ZuMpdRDCEoTlO+dAPKJIBkdmqL9XrcErVGLzttZ4QgvlIFS2FEbz7ytGdfjpL25u
e+/p2Db8ibwcSbNvjxc3cgNy3c5IynoPVSUY2v8f8fO/JAZilTuvC6a6jrIuYfXx
UHzbph2f0045++hAPm40NXq3rqxwOmAlaXVLRCaQPr+GIyTUPH8h/Osbo3Yix7vl
kuDqQQRnq/k7WZEH+7ZSjORk2bQpI61yY7bejqoMMxJWjIFTrmhHc4Qk184Rq1p1
9q7rdCXWyz79pB2H/QueQXCLuo4bFuTn1ioVrtupCpm5MXm67qaDmhEZNIh/5zjw
6nGbjXgUY+UQgYkKMsbf6JP7a4C04aKcJMbXGHIcb4OnkB0KPX8Hzz2nhhTqqpUP
dqcZD6I4r+VHukLnITPukD7lX+ZWeayZzUYpUC1M/d4IbnS1EMycje33nqDyhWuw
BnDSY8MaGdZhUbQAGJ/1oIJMIdGRo1pIWe7FSSSeojhIDKqXCAG17yqygFa3Na9T
aOAGma+UH0LaGEk3GUZyGwaTVZSRz+iKqf4ZQUmyhe6YFS9gvn/gm0AtW5inDozx
9oPUF4JZaPem4y5wNilffVMSiapWEsASaEjIrf9AbS+fEoL3BlwvwzfgPRT8xQ9z
wDCRmROCDZuiMVwfRkVD1YGUJl1uCzgFBPlUEDtAI0GfApLlj52dzDUPVHlKnDJr
6jjeftSMW3hVFWlB35Wvs/jGOIW3PgQ7SYVqgNUwe1AdoR8LyHre5jmRmsTLLaT/
Wdws/bAZheadiHqp78Ne4+ph2iGVeM99dhgI+Xzy48liekT7Smr8QZZwKyE3WrTf
XlrLy3wph4NVhSbnHc/bmfYoqEehdOs590MAMkN+md+79DyHwvA0OKooGVPJDPGy
95qgyIDgA1xZUXVoXgqpzvytMv6NuyG/dmn0J3FxsHA3dMilHh05rkZIkwBm5GcH
/340RsC2MygX6TQyoTMz3MG7UiQCHIbcheNbnSZUu4StdeGC6lqQ3FKLkJGtc4hc
CiZsLGXfS31oPwkuCMKceEn4B/Ct0e7kG3OUgD71KCGhyotcwvXODkUMgbjNJAz4
o8UgIIBNI2pndxTV/CHSkuAYog6RNHLm4RBJ2SjEPqTLVUvUaGcodGOy8pM2vG8P
wMJq//xv5lKBVWcCdFClCebs5jvHYB42MKOQby1TeR+qffkF9ZDev6j6Qw0zUh9K
YbD/kTmJZA9AsoQFxPKp+MJWGbO0z47oYe7afALyasWNNV54ykwE6gismzdJgoE3
CU6JUP10ITvRMDtjbveIV0mHnMh36mMoij7o7l1PJIiMz367pPQRsTSBFir1e9X4
NnXQXhm1heKlW7iMpo+Na6wd/1Hhgy67lw4hwoo+7F5xElmeOqAVwtpiilQCFjIu
II9ak01x6WrWTi0J/8o04pu8y/RM3kWzNsBsT9RZmzgP+KJyaQQdiztUrpwOoK9F
+uXoc/0Tayi3kKCWRrcdnZ3AhcrqISrJjRdofwn6Of7L1ZSTK6wC89DUzdGncDay
rdTfsB8V9M8FyxxyF1o6+oS8j5lFESF3V1yr4USAuGygsYujhAcv29aWLIz2GmdV
yvduA4zDGW1YRSbPr6zpQ0DHG64xv8rFbvsxX9GUZwjxtxc4ddfp7p6cJsjagKcE
+6qyveGigfNBl5MMx8sieMjlp6Llv6OAiOzOHVPZKfmxsYdF+34blr2qCefdTpZp
JHON+HYjbIEzok1BMulCdFSogMBMHmypm5hEKDKlFf1GVRjgdYCqWksJCukGUM2R
sCUCs5waA94zVw6GhYkFr6986QWgjysDjVSjGmCnWdC9wtaVYG3BnGpkmbeQi1Gr
igMKlabPfYhLF7TAveGilr8CK50QqQKy3y2JoFGrwrI/ngMWAckVZeOIRvPPIeM6
Xcm+11+bmGhE2uQMogAfjP6Y+69D6A+9y0QpP/2dUn0H8SJ0IYRMSzZ5LijNi9hA
EJ8JFQ0RY59GUtMOdKDEk9yIvB9bGIysVbyL0SuvxLjIFDV/m2xnChjhw8KlU8Wj
K9zpCNbZK41vFPNlbeK+PFBesbhbjntdCOaGiyFBZVhweMUh68LYFUdFXCnhlRen
CABtSB25GWL2E0UmH1KVqeboZSk9zFrt1iW/YjOfplUo6J666QEZGf53Fc0RhZ1y
8v0EsJ+A94Cy39sBrCjXAq4NLHxr8yQ+a4lpJucZXtBNFH1pKtzIGaz3YmtDffCG
6H+FkQ7u/vwVIbB9+ug2CeD5GudX6FvvEeNGLrmHE+/Y1vTja+rLw+tJV6aja7gQ
ax8Gme9zIUSUG8FRFkRZHnZQ+PyV4ZHKZXMkMqV87abj+kW4SpSik/x3LiXcz487
LcPz+vE8MMmdSaH8VrciK/sr9Q+IUtE28vI2sAQ7MQCkazLi8AQ35SpBN4z3UmkR
PX5HBk8yBHeWCtFvkByHMeDJIgJIUkT6fBBJ9MszPJFz8Dumve/r8uroiVYoftWj
bvH4YDmSr5vaiQPiGWE/KZu5brgP1ljltY8Qg6E7/qxmSCYMrJzEglOSuP77a8Op
steQQeMC/825aiVr1ZAiZVrD8S83PJWNubtqSLdlPl+KRsRqFJ3vy7O9A82Y0IZj
CVypKa9raCa01TQiIEn5nlkr2FV/jqu4sYMGqFRvpxUhSJFNabxfw6ayOXQVZItV
5zVw38xRkIpMaCx8Lov6DlOUO2rSpQefODSIu0m0auXLDNgpButzpLmk+JI2WEMo
CNaMcKz/luRiQCi7gM1hdSLlWO6xA6zgBZXzKaA7u3SJwwi+ZJAN263nUWK9TTje
oGe5+xpzt1rGfW/RLDmoiee/DCvpMc527FqJ94/6opDoHUJNODsZ66mvRUQPF3g9
0B5cqd7uEdOiHKGffX745F88yN+f0nfdy0UMLy7ndtTZ69cgkYhothKoDWkJQSgK
hgqGK6i7tVViEkBBj0vaWF4kSORQD52h4Ty2fVqfxSVb432u95X83GDOpZKka+P/
vbpHzcZ4sjVe3baRu0XfkFXo0qBUwsPyYdmicfdFeYshRiU6cl6MmMM+vLOBdBK1
G6BOYJV/rN00pJiIMkyPgtSc7TUhZLhHODHKZsj7MBL8ii6AT4xYWr4Hl0+z5YBm
Awz5++aggBQRMcNauXV1F2RvdL+pG/RAdx+drL7kpP1k3RZwAsQpi814x65vDC/+
sDlMjEhFMNLQEZzXrPKt8NaAy/1aQql3qfGRhl3XqoLNvdzD5iK0ihUjH0ZMSxy4
R5g0nlvDuyQkyzYwk63MtHre0hI0Vp5Avr09ywhOoTWnqOSNDvZw2ZVlNlTGRG4v
xXAQhBDeMk0wIuxdJzE6heyRaCimrO/P8ZpjLffWIfBq3D53/e5FLL5mw4KgYgFQ
tjqSxjHy+OFBYWwvbjaORWE6KuuzoFywIDKnCXdbzsJASqkqO2zpopMnJynO4pff
WYlFl6WOy6norl5+izVEsntIjfETJU/eH7NPUkISTMy29nQbnD0+ZH6MHuEk6Tn8
hQl8dpsKRPTZheWzK9C+c/unX7i804FUkiWnyQjoBeqeQKcevWMwhY94ccFt8U/m
twVFUOe4/fyg88ArjTOxU40sVzfgUxN/behYSO05ExDlVhKy5iDV33d3r6OgDvC3
e2gM8FDx3+XRjFiUz7JAJMjQZCb9sjSkCICC7nOGTnBE6O8subjEzJsP9tb0+oh9
PuK0yt5VqQw9838rc1bXXwC0y6untli9c3jhR+gLA9/ymkmq4F3XYhPDsW0vSveg
AQxCLPUk2QG7/E68hH8iTcFDg2LFZ9A9G0+eU52n3GS1gavxNj49GygfFlJVnR6j
eQGhOMbHa0YVBezn1/O3UWO1mUI0ZiXcN921kEBicpZ4rUcNpRIENvz5tiCWIhY6
qEjh7keCOYndeqlOgng2y7VWXpn94fK3FsNxEbKjt1CCPGiBn9ax8RLSIGP4QiSE
VDWteLR5Zy0+jJOiD8KFNoiPsYvLK6I1k3dKiihmHGs9zdL7QDxzeqYu/Lk1N+uv
BMW3GdwFfoHHQS5TSWnJmKzQCSMQwuB4UVZGhQohpq2IsaMDlcU3oGYg0ZJ6IkXO
m5nmrEp70csjnaQ4DYqWvCZYXox7aSiZ6cSl7jyPTD7wZ09zIxs7vt2UKBY4tKfW
52rOxO/Je0/16rYmaEFa1EKx3F0zMUv+iQaS+Dq1LSUbmeu4CJY8JhRNSCPkoa7M
pQFPxh4PHZxk0OfYTSLD9kFJavMaMUmuc1jKJWdy8mxfljKyyiKTJP2R908+F0OY
LT0fhFtcHimAqBkvu58vG9Jo6U/McyjSUrIir4ZlPki70cQ2BrtmmT25AGcPYyuz
r60N+Rj/q3PGWPfPf5H4+Zzqp0FqhMjv32bJK17140h8eXdemsxgwF8u+x7fkvWM
YCWHm2ZIz0+DlVHLxji3t1uxHWPVFLkSwyVzTPhRFx/Araxd36Y3fTwv8lYvSTiA
ImxzgdElKV+o6+NTR+Kfp/nNaKF0mBGsNuNUvJnf6hBnZjHI9WF1gTyB+tjqfo+n
yddvXKTEM1bayRdgSOtJ1P/YADpxxUgnSaK98OnxL+itFxgMC0ynkzYZGRzIQ2KR
bI+wQqvYfd0XhycT+QNuniQkCdrrfopJvGZo2iNFL4CIp9qdBNTC5um7uOzlezie
+uvUMIta/Frw0DIDwgLzLEitWmFPjklyu9OQj1cFrnSNEhgDKmnO8JXGqdaOHhCa
fmLs6I7ydikxu+8tZZHWOhK2LFlTZBjSB+BKPgX0eNv5PUpRHrpX6Jnl/nZeAFon
zp8uqpc82afysy7iZI9Q8b7BmC0K8wa0E2XHUcRG372FAfqcdJbzCpzzPWgbXpyq
JdqZ5pdYUMqfWq9Dh1EA03zen2gVCPMPB2xDKvpSJJjO/FeSTmkdQVL0YatNVFFK
S2lb9OR2dumQs8o/x5d8hQF5E0tLYPJ8RII/hmD43/s9sJQbuLoGur95B2TXezYy
UMKQrubH1HyHCQfvCwSpU5xM54UWyl/2bVkDAp0q7XN8UBxyU0dancoefzPFUQk1
7q5JsMyC/LPAXJ6BB1l33RRgzCF6512/egNtyPU/TBedzoBDHCb5UL5Rr0vARLBQ
9dnnXf+BHswvCm/5lssHkh0/V5R9yq9qfwtWd6yoFfC8ZC3m95Szh2Cw8UDt9QDw
Do19x3q9GGvDZV0DFxUdvXnl/qP2AxzuOuGL2VlC6Ko9zLQQEcZsUOShg+pOzpdO
BwkU2/98jN1kzio9AXm6cOiitMUUfSw2Hs1m+3ktUJ8f//O4MKpb4Ur0IrcbCIP2
/DvCVk9U3SUl10LaWfB9haesB85tiQRmXLbUCimLzJpgV1QOiQfAdQx1Z3P4Lvc7
EyTEsidN/WES9gV/6WHlwPwkVj8UKU5z32LlsQdUW0UNLKjs1mbNKssOvj1rnpiF
Tpdme8IyAdUvYRn8P+XkuLkm6G8RzYodWfB/ObsilnaAywPx+pLMm6TVcmYd0ejt
P9s4aagfZJaeExnc0toYjOJV6WBbfdeFBI5wKtFtRt2wAZ2jSYptaqScaBzr4JC5
Os+B19/mw3SWAJ/nwIxLki1AIMnA15opwL01HHh1zcO6YWqE3LWwuPM/+dh1L/eT
fPf+KrNfbjmw2ooRaOBNEZXgP7qxeV1cB3OAMLcma5sCV33xfCI5ucGuihp+qmCZ
0iLv4wBVdoE8EdxHOTDpgDaDu5Cz/osfls8D6GruwzIQ7tns0X6FGjjF9QCEVbMY
E5CZJS7CgDei/K0q6RusbQqaxCi4fvSICEExP2DZX5ZgPb1reFmOw4mTHopI9jWz
Yl/oYdDIFBwqXMSOvqhZDp96Iz8T2KPWnrqDCsDErCgyu1xDD9AHXIRjHo/R1UZ3
imsdLl7NH/+ZlCLf/ZyWKQ1NFRP0+ntv25M9HLfFZ6990Wj1IY4xVfMdnCo8qz66
8WW429MXNEAyAQ+xy/osnDW20p9+l6tJduLE6SmLFPAddK+U/7oTDkRckSkmEIdl
h8qMHpGsIvkawVNWJW2KekU4/c5tRP+4i/IH3pPkNKRu+jIkv92EUgJR96Qg3lkn
xLU7oz3nWotY3ysW3KrAroZAyJoyZGzVeC8FYMwQwWdoe3aJGQKZwfvCwytq+uE5
rPVm6PO4YBZwmVSNWgQ/oHsybfP5kxMhcRhFAP2NKHTwKunOYjfl+42kChwIUTro
dmyZjbdeqTHvx2zHQ0UHR8kAUQXaL0LuncXfFe8pSYyFKK6RF+dhVcUm1GK7TVlu
GU7ehlfaMkRCMpoQrTltur8Fm7CLreE7diiLf5FS8BLHW+um3zZmKCBxSolVRxRy
Vpi81Vefwwp0ZZlGH1A8Zb5ZG+Widxj5M1xlNub6MU+Pw43z1e0INwSyTmx6CZij
yy4gABGENcl+X4kHCmW0egP/fungdXwYWnb9ZMSoTXqA9pqRf/f31Ce3c0eTBcTG
Mkc2Eg12C/HlWQi5v56MKGaUizcJZPWr7fXVxG7eANzUkj+TOZi0KB6N/SyQ6CFr
evlX4G/xWz2XEvOjcMCaz2RGC2jVzJnKhBIaZ5ouSSb+a+3EYOjqu1oaiPqlA/bL
J5U5uva2w/Ze37o4hKzoVSAKYBOnMByfHqZbAQHO8QLpoFrpAKebFtPG2Sth5/hD
aZvvqhrDfQCa8ij+kB5BumrjolAmD8JzV+mnMiZd4I6qXPmyLh4JXwv6x3oCO7QK
DEEhjYf6g0lSSdUAusB10wpixC6i3LuPrCyhSOE+WVQOMLbCxeMmD0IgXFTXFJ6c
ATyG4UkP8QYtJHbEGjGE+wYk550eq7q/1+f9NOypSXrVk4MNb5huji+uDe/XH6CG
6eEWoE17oyn74XSHFjWbQJXjp2SLNiy1+rz3QjXb+PSf5XA5K7W22DWVxQdbP8P/
M1IPepBggHfNwmfkJmNrPkauZuW/5MxC70+iftTbxbi5VgJP16Xu6z0bMjNbzkhg
EM9NxRT6zkjYKL7uOVvUj6vEZ6icPJsaHHEgJ1Tl7SRF9PmixJG0oFMMTIqkF7GV
COkSgAiaOq0Wa5dSDtQ8s1k2jn0Ahd+s38EtXIim8LkvNuXxS1WuPJLWCee4e0rp
ZdDTlgnQdOFb5OXAW15+xy1rWjPUGgcelRkXsTE7W/0cp03JWALp35RbR+VJsjzq
QhCCYjwseV0zRIXBwwElBzOXv+3MVq3ief4ZaIyvZBaAcoTES+QYPjLVlSsQjOgu
DwdZTy8+EjOrKy4wQ5UI43vlO5Uyr1zPgK1/pW+6emC9ZjxBKoDaWxzPWrRUZW2V
FypT+WymuMY3B19nXfrseKkPxTt2jRsq/Z6C/gatxe6j2JSbAi2UV8TK2sinfUbN
YDl+e538tjZgiv0JewVRzXAbWbvdYbGpGpdidxaGzNnW1S/8arCYFOiBrW+lw+vt
JWFWWoU7wIWJMcgoFXT8gedN9x8Jf8+VpjbGq+PtyI/IwHInd3wxdYwafcDLaMdD
xh1Lq5V0NpGwNrZ6arwMkXog/XBr/PGPjPYk8yNG6GJtvGbe71kElzD3iWPK4AQE
cqO7VZgP61DuRcaFwiT/F8OXWjBwfootBknLOCRmlCRb8Xm4Dfs674+0WTWt7iqW
z+vgXtkZG13oPF3nFrpXaYrb9uNKWZplirkuPQpSVNfA321zoNLV/4AwWSWdQ4h2
fP94DpvLEPyY0PkSEYfqSn0zjQZsJkz1GP8ZsPCVetWl4Fn4vd5Ybrg7ExUeDrye
3K+MN/m18su84V3Qe88ErZ2jN57QwCDLj2Eczgn3gdLcmkT0LCSLhf0TcHzsFkpN
EavZdsMI+r+ayAfBUzenH+lO+d0xWjrMGsG2hq3Eik7tXlzHXijcJScDKGQSXKFn
uqDKV3PsH9dlkE0sbjScaWZrQuW1HGzBV2Xjb6i5ZF0+6ENUmZNu7IpyMp3ROqyI
MsELQv7Knw49n7YFt/dykEV32ZtqlXRbCzpC19HsL0zJQ7TJ2wH0HkoF/EbZW70T
rder4Hy/2F2v56fyNsI4sWfkZoWMD6jAdVGs12FXX0hCPiHjkCMDZjGZQZRaXpGe
kqxH79S+BK4Zptf1NSTJxIdwxjoe9Hi+JpeTnv3FWZQsDzY1hxUDPdr8CKcKefMR
DvWkoTAz/1xwbCv9Jb2I46e7PciRPB2VG1OwPTcW7CD5PFkvse9X4BMQlJQJiLzR
sJJpfT09HDcic+bl8uv/ketFLk1nb2UwUITSYOQxNz6F491cRQ2HRzTDOmFV7zki
0dOA6SGkyRtgM7KGMX6fmnRQScXWUV9sLNqcERnD6qm0tAEHH4L16fKx7oRW89NX
LpWIQq+/Dod0K86kFsgjYcGK+kOFqhB3fPelbeh1AtdCkSqwDJDm0OvrQWsGWH7J
nXGP/JQ9eB4FMht690obnBNXYzCowxMnCKZyiwerf5Kau+fFwEXexV7pvyCnKe10
IkrLaa+Ce0JGxSu9OFm9Ai3bctUxaA7YbqnMXguHifHghHEcXOX8JIkEB10m/Ywi
oWMnYw7+TALDU9/Hj46kOuM4yxdJBf9JvB89n/Dfhdx1G8OuUsN0k2NcxMLXkaAy
yJ53fVrfJRLhwyE7xdo1z1VxbPq8vwrZ/mtIhXmLKl+FK6I5VfSwIFGLEPdK0qf4
YwrvbYiHwzEuB/6L4YgBakLVLmz2YPxGL6hxtUg81r96JZYau1LIfNf5vSo9NlHp
RY7npGG4nF+rxEusdnl+oftUDDOudRavYKYyMW+GFpqJXpyFQFfFC8Nd8+pdGRTs
3u4fu6AERqki92PzZ3Fs0dv6c8G9rEm85/urGBTCiSLcl8x23ODptQimmO08gpFX
1DCVkiD4sghSFWI1wFiaqcjVxQdhH3ldPBVINezWIZfPzrGiUQAZ5C17eD8US8yq
NW0eRClOm6ma16hO2L/upc3SMSL5Zz1kHLKfsQLYtGlQ5Pqo0rVhsTLWOAXHJq8P
Mvb/gebfGoAsuQe6XwDRZqJD6JvUj2RKQIUYdYaJVkx9QhIICoNlkaIK3Hc/aDqC
WTM4c8dM1dM3Ozs9WxGyDMvys2eqw1oOrv/pSqqQiKp7UyM8o0I7ttsnYWYxQQH3
Cvcqz246az09UNH8vRePveUb/x5tv0XzofeTynj5BHiX76+lciRgvUSKRN8H83CY
4bHuS0rQ6DGkGM3l2UUI1/SHrobM+2FbW5cquVfV1ELNuF+/1oPZCarKA34/yLLD
GSEGSZRZi1ucretO2gDUDMnRSBhkLD6YNLHeLoGd5liVs4yHumLjOxfModBAK8Cn
G+hfh+a78RPoMAb/Lj4UkT+Z6KWLhr/dOeFYHRkKUDWwQixsBDaqDUMrb8kKxu0D
Zra8lToVo017gp5Tc3uPszQtno+VUGbIW1QacH7Z7gt6oYpaBZCMfSdcAz9Pli/2
Yy1S/RCToB5nBnL1Lw+4HRbjlMP1J+ROsriyfgIX2WgJuCdL7MrBKV6zs2XVaWI1
5536Rg450VOnS+NBJVA2JE/XvzCzcMElv/Bstr3YIFD8PStUuI9VyFViXt5fo71y
T8gwE4RmDTb6QWRQzJ1dKjh6wYzwJQw0SeRumF5VhHfgFex50Uhu7LlVFgWQWULb
1DZ+lrlVBS2UVQgrjLRsXrZA50klyVQwMm2pNJI46h26kxvzmNBftOPku84hsQ7E
sLpiFDqAXsGr6DEFdPtqECy16sB556eJliwyvDeBIWBlq49FyvuEuZ4vlKsjnqbQ
RER/qOkiAVq9EJTCrkT2bLY2FkR0E8F8q8c0/t9vf0S04OHdAWoK80a9x1rtj8L8
PVOmlAjOJxBaYvTWF/2NTwarp2hwR1v2d15kSdZAQQxJwFKdZdNt2Uogc9zlxlHS
SE+S6UdRfZo4PQSxz1iHTEMhYK10A9/jjLpr01DqfTaumkcUYyYsZigVjhWicTVa
DAqm4NZZKbDgRLn/r9zYOqG0K9s9FoUqr1DMzhexd/hErotv+6ZWauOeHgNibKYx
+sOx95Ed2Ho5ifC+ydvmqEJ82r6HNHhCSprynFkDfLhJAlfCW1EFm/kN1UHIpFwQ
xzmALLp1knrb8wNOKyI2squz8d5Yx5zSKjFqUJvLt0rRAxuwIcl3a2OJ5G20u2eV
w4ZBFZB1Aitii2U+o8J/R1ADyf1NAaDZxWKPtAiy613JqvGFUtxPav1MaAYv4T8P
D2BRewFEB6qzGqDGNz/k17GRSOAym7l6VphHe2AAtvMqs2Hp05ipInM4MlaaTvnZ
jaPuF77MQckAeir7/BjutsYVcQ5PRETmj2c6Df1qjJ5k6KfwPDUrul9VPwf1Pgha
4K0CRZACHZWRj2dnMOPrVt2usi8BblIlH/qhc9jc6lMh8N8iB3Fyv+NcaxoErThI
cQ35QXS2gBYNfDdrSH/quCV9S3ISdf86754crx+jXs26fcmxWyV6viC49anLKN7h
KqOq6LSnthmzkmI/f70DIYP9qvH+GJdKE424yoqKhfgPHjfF0x2ke/p6ZeTyz6JZ
5p1y1HOLSc8X52ogMs/hjfPctPOoOKYjKsaB8VfAGY+C3YoRwdtC2WczERt/3xdU
TeHZUdlJ95MOdDSmoNg+rkTMY4qwbt4ikxp9HWe5OeCcn5/2meuVcyAHNHUucybZ
i0AkwS1aO58ZVL45UT8JfMSy7O1NTVT3iP0q5AQfzK7lATw3RZO0MvQKhOjNwU9B
+5s2Oeye1/37D9eVhTcTOBMUlETsjdHtZpPb+KwHhHM0fm5SeKfRrjYr0wHcEHTK
5+tc1DsKxFIjfFpUuVx6kFfMxkSLXvVjDz+0BIqWQGyOq7SLoW7Z7MLXnQ+ANSkA
SNZrvOytTb0FpNyVYDbNAjdOyRBrch1dWFkVkhsmWE72vRYdJJ4Bn5rixImgytNf
9c99Tj9RP7BwjgsMs1GSCYsNJKINf5ZdE6f1hbSJha9AINuUOXUb+qw2+OuP3Pvg
6v8RqoM8iGGE+qfiFOxQFJ5/xkcHPjhrY6JiJzytfQ3/TNqdJJueh+T841d2chHy
B47PEqVt7sZQuYtEqRPA6A46R/MD/nTMhI2eM7JbQySUTUJ+Q/7s2xFzyEJ5+uBp
uUJqYtRRGJRdjlnwqq6dhcWu9pyM2V1aP0V8MRidTHUiF5JrH7HqYm59HnYr3PUo
NyPPL3qfj//LkgxsJp81PQv8SCPUS1NwcrPkjgB9B3FrjVFBi2e0IqKVlgQbpUy5
XQ1zSsgD2BWI8phgYfY1EV56fFyrLYnXZFG9XRV3sFs1HrOipgBPGZiHugj+meU5
41GN2G3Nzf9B4gUTU09mMRJmQ6IZX2q/Zdxk4N6mw/tZMlN0UeXYBA4ei+3eKOkz
4gf6KuYZCtNjLgjKdsSdb/vpFnJG7R875zszB2jpTPzH/+tfaIorgMPqZtvLrVJl
fv32+wUmgNEf9m3cGXsnjppNhwDnWjCM/7NDjaFC6jh8+biAIjipyW3g0D/s8aqj
ecsJ/KtE8edzUIYVfzl0xaqRBTcXVJ5QWIBpTK4H0HtXt6eYrzyEV5yAjDIZn5Mj
gScNaJpE+qQ+pT9CesNMYSNVWPFStLi9A+akPGCjxaW+LoHL/jyS7cVuiXY82hOr
HXPDEUdphV2/+f/oDBZKizyCW1Hldm62EZe0mWdVCBaGD0v9SQIjb+zJMh1GkF+O
ByYFK0cxebNLmdrhl+LDVYuQSchycqxyTctF1E4nRit1esYALzZ1fRq/1bNQuv2l
xs7/CrncIxvXWmWodaevS4sWo71Rn6XtY+sQxq7PgqIH4UEMCa/xUPTwJTG/a9bc
5wUx8EyOX7xnmzvM0ItK9aavjdPXBvhAMgzGJ82FrpBR2BZXmyP1tfe3RqwatbBT
7gy8efO3ludog8s1HbqNEid9cQNQC5bpQh659kPciuy++/yrZYOJX3iNjbYhpSHk
8uGNcmC17ayVxDk+dYvvYWc+iz2qRHnCmcg4nKR8Cg0ipzo+AGVU4NUk6mJyiv/J
mHDOJRZYi7RR58EEOqzHTuiIwpIv/uUh8y+lKa41oauXoQ8+0x4nO46uBHg9xW7Z
KIQjBdYxlHZekLw9RlDy0XvTN1doqHVFtNqQeQi9WiItSxxCsbvXw9NvPXtYq0HH
/+0yZRSVSJ2/ugms+xZZaqV15CFWfNks2Q1cmo9Fn8d8mP5UwpNIawNBXygcRPIa
z4yy3eHFbcCa3h7A/HlOdbBFx4q6DxuU56nzbFeJSKgBWqriOq+TvM/aT9HwtVPa
XzdIFpnP17+tgwcXmMhkZNsi/PKivzOdnm9wvOoDLOojRLgzRkjOH+2NqZVmpT0o
57N/mMkYGYWfJ5KHbbILG28zzLbkLHEz1jK3j5rdvugJOZGcLhdwhkQAKF5tc3Q7
Kv8GTEtFcrzWZCTdTdpBHNb4gsls62a15xDBO6OaqSUSI58I2tLFUPvGFHb+mSW4
mmbeUGrYQ/3nKSKqIEojX/U6JPYxl7aGZIDHtP0X4m38S72J6TBx/dsFqeljh2Ou
fczmQXcWOVJXP9hlpEpLlcUv+0HI8Dq3gzxgh6YnAdizv0OcttsDf9jX4U6Ey1K7
HTG7KiqlAdoIW2wH2c0YnizazfIvy5wg+puaG5/Jz2ku0zzHUmcrEExbTC8+ro1q
VLuHP9YI61DFRbSQ3BnXG+leQ6icXomsN9I0MxovOcEgBR173f7LKpLAwtNiWXbp
QLDt6W7GcMMSKws9MKr1b/lG3rEjONtgjx8+tAAEU2uHmuntYbM6+ZzWUoGe1zYm
jdM6CCNwNKJvN9UwSHWN5FPmDmESWxdm3rH7VtzThZWXGa6bhdWFLqsH2OdJb8RK
X6XD0EeNwENbrpdiXYwuLipZJJ9Q6XvbE6qQ3EHQS4NYZK3LOPLzb6axn6ZLkPXt
D7ElLLeyMZzxBctdZvxxDQdSQ2mkDUNuGaP+zsCmz4jZJBGXqX102Iiy9Mh7VzcK
Eie7hbyeGsLVvE6olSni1a1KQAegtTAp+cJBygXeVDslGRtYi60ysBZmK70Wxtyk
H4aIMO2gN0RwNyKp2Wti++DAtlzB5WvD0/uI4Ccioq8qR/9auTGLbpoMWeI7MtfJ
5I+fnTURZHhUNlYpyCtDaPoxRFiwliUjkIVDHtAeIdm1hA8SLu//fcGEI6l8HzBD
8H2hIa4W1JwyzTTnZI0Ic8xGayLBnDkyw805rAsV4gjOHBGGUC2l3/2pqRsgKkSq
jQuZJ+Il25cs7gRDVr7G1WRA/N4FLovWHbOly2HDi3RMeJQsFPLwzcIsDav2LGja
dMrSYArpzzMjMMUaqJT+ZxvCdx1qkBQ2/OVeeEEiTuKkbDmA7d1fW8o5W91chowu
JVty1nGw1DeuBA510c0LV4jjbkpFm0Eilx/SOaWTLB7nbizY9KkhmEE28ahD4q9C
UOj1bPyzCsKXvaRcdahBZvJTPbyG2J5mebBC0Wg/SRhfdzXMJHh5ECj76zzQBT9D
vmOr5EZmj+/IN4/fsjXR9KI0YrR9WV0oBkGUAHT663dvP1aIqRSYl2T1wF2UNfyM
9h4aktKaKdDKdihR4r1DX8m5x9m4suSFSWUMPnGL6uoQm+7LUQaC3uQey4oFhStS
GYcQ2POxaNittdFlWTZquXRsuOUkNdVsfbUDHnT0YVbPlBXf0yRv76W3j2cW830f
IG3h2j2llEmDYa1jz63C2C8rg7o4utiSQfLfm16ula3oTiqlBFDt9T4LLQjrgIWN
kushgFkwbArSPzPzUsCz324MGzdwywzaIYUkJAT69IAd3KOYJIqQ26LWBbI6/ZNV
wDre9ZCGI5uAMzdLPHyh1zJUa7jvjBbawopRW8GUpQYnCCJAQRtZlx0ANiUqM04c
bbJPaVp6dP3IP6ji/kqk4kEQZ2Sw/RWUAqQzNvzLqa8Qgr26hXbjp69tF63UkKOR
WBip98YiEwIufgVLECJ+FNERDGjjPnCGoBuF53haNhC85w9NI0RoOSTu1B2foDBf
9sLToTqKNhcw8ayjXJiZN2VcsPXSBQiaSIFw+bJnzFmR27XSzMlcx5xgfD6eaz5A
OqM7zBOwLeatG6u1hIb1dXsIb3joIRe9AblBVafBTF5b5/VeI8rx9gG5geEd2qan
5OPQ2WTMJvqpmSelbZn12Y7mSByGHwUllANqukHpgoT9cYymyRELmtTVl2bWgIDW
ndfaBBFDmHXfK4rmVuL4DyAiBUISWZiA+mVWz3QEesTY90CRPaFIzrFISzVArlvx
rqKmiwAf+TA6qnYL4yqCVZL3+KzE6woJyyGsaOBw1s3bFjbYpwmGVD+nVsIDMYIR
FKmzDIyIsf3T0YUA4w1Pj3jMcYg51ZscbgDd4Qip73v7Rxb8b5SFQZNPtruUtREo
dNiyqS/2VPbdS1wMoW2cTx6l8erWefilFXoLg8TjUh1+5o92JuXMsiBIgLchBt+K
eFuVJkFz9FGnrlTGxr2viQL4qfOxqacpRkk7mUD8Mkhw3wBwhSGqKprJORYOpG+h
dXoyCGN/4H/xJ51r7ZdkE3rWHgJSQK8Bq8CxqJZGqCROIQwrDvcoBXOnAtMkuAM7
3r6/XmH38ZgTHS3XA1wzDC39paTDwciHSzwjMQqTuw6tsY5mvi004In+R4uu2yOw
X1Abt0xBqiFOGQFIZy85QIGaFWzCAbkAQRYgrw3By+DI9ZUp3BT9D88Q2bt1LKaf
tmXCvF9xTGFRLkPE4URknF0NFuhcQ6dsJ2tOsW9XgNynyK1+mFlnJOr3XTlCvI+u
q0dfUsQU18aNRVy5uJGkfWoML6fUKXIhT4GpxATf7xiolgLDNKTFfwb7p8GkHXHZ
umk5fmT9Bm29tdE/gl82InZk8sJeoNS81NF3Dy9k42FgLXl41LqgWhJwQgDdKbd1
m1CrC1dXn5IWXDAP258lQwvr0xMNyj/l0eR05WW731xm2aSr+YHMLQ60WqkXUB4D
cxdqd45YVF5fQ1KCcJs2nrbKNJ4bx2XZCq0utgLomYDVD9Z7pyPSwv7RyLfAwzKw
pS+MS78H73gb27PpjC2yidvoP4VHrAa7ra933te4jJUtuXmXufRdRfrWFWezxRZh
5M1mosSE9YprbTIDgU+JDqJcTAkjtPRAxzOwxaI6hXKssnGEEYkkYW/SdviRiUd5
s9fKBgr3yGo2X0wJ1Kqm4L7w1DnyINMNbUx7pqPsf+Bzt0IEhxvhjn5AZAJh6boy
FW1w8nbVTB+JOu/ncpm7fduGSv9ppyv4v9hfL9aT4Z9hz4keveozF59TtB1bkM9i
ySc4ihDX77mvRYIfsnKxNIvykJgoFAIKH8K0I5Os6CTylrP2ARad1eFdNmCMvCK2
3JKBSZAtu0+kC4rk//7vtjlTaPnmYTGcyZOoyt+E5SvpnTdRJNn77yci76uMsDHv
5hvGTeQXuCqJnorTPDXLvwCyrAf1h+ketXWnpp8MPkcj0d5edloqDBAIMokuBXYs
k7IdLGwMcaYXH/JQ2dVcxNCGUZgLcIl2Z864t87O8pBbiky8KM2WYVo1ioPxrzMH
ycbB5hpZJ2GDYofPeRrVxf7IzbB1gNK7Wf2hx247OM6v9MbarButCq2ljh9ZGVux
hGMrjzZ02s3KHlLlZvwfzgNYG6YjEoKEd28jB3q8x5wZTb3Hu3SHcmXCDvXQDWDh
LBSg+6thg3bF1GHok0uKg2EJiESFChReIYpwRnS0Nk8BtTHxoOf9U/S1zA65Fx8c
wUy/Bki2hznMjmvH2696uwwaK5MotFFCdTpPG0urSOlfThQl+mNfCIKsyJ6P7hHq
4jXRyEciNgqsNFQ3fDt7lPdkJiaA6djAw2rQQcBy38StBpjSOZ1I/ctfC134MQGS
mJ3lhzX5QnWIYgJrDIHR5cG6aEZmxk0UvZzws8OVo7zh5fY6+dSyOj1pXX5TT4+m
Av2xOD3Atq18lzwdaIXAxa3jL/0sr3Lj7BNl+awmSOx8GDOTNk7AGF/sBWfLSdXS
zkamquESIX2qWeRibgXvI3uLAHk4x4Z7kIq4ok8OgrJPMi4eUyjvhRLG/I8UU4QG
ho2e47xEUs0oPDsl3GLXS24GbPq3og70kTBqTEwFJJJSuEQVgkERfV3NXrtB6XUD
wajFB81CiLxPIwEKPHBJ2VrCeVqjS31Ibxne4Dnz0j/2WhR/gJ/r13UcE6fBG2MG
CaCCSLTbzFP2ENWbyFGLRKNhpFfj+0Pt9kxhwZA7otIemMl++Ex4vCAGF/GqG9T7
nMqOAwhGu7hPQcE1PGoghfJ+hiM32Gjbw5napciq5ayaZjZg3G83aoyiIf23dIli
ap2T0Sr7NqSYdycyEGoZZcXtS3fPcePdkwPTgDYcc+/22/9e9zw1VANsHNsgsX7t
gKernUUncAV5iynHoc+aCjxLhqyi8X8l5qMEDdwmF4F6CEII7+tWUvdFjDZPJCYA
lOXMsuPvxZmik1CBE/BRulPIZ+Kdzk0dNhDdq9vgYSwHJ8vmjRhjjS1GVyDCH83Y
XtDEl9tJrq37U0Qj+20RS5UAS2dR8MqIgE7sosTIi+sIXsMW56clcL0tugL4KPj4
odqfA5L95gBk4SX3wWuoQxOSGm4IigXIBcMoTIJIEAyZONKBvxMBBGtjoJ6p0rhW
mHVYq5NJX1sOEh10YUEHz6y7QaVDoxcrejZPggjgY9w5J1w6HlawNU5qTwClefCu
0WXBjzd6l2Wctz2aSfBXTCfmbj9ELj3R0w9MMVf6/BJc30QWU488gwqcHQ1Ug3Lc
zkSamnqAZb4mEY7xNzie0mKEMfWharVxh7dKsBjtNldDWuVw+4txrdtn+XTsWsMS
H0iovHl1Di+3/Qqc1rDx8i5WvAghp6oF2VVMeZ72X0o1RkdmaVJ3br22t3pf8aj7
uFh7k+hjhOFsqGdHc2gJDAGbfcc65P8h4AZquLgkSTQGuCL8A9uc8Qi53XKv1wSY
Ko/B5H0DabZTqak1zGLc/BD1XOcL96Z+f2zmZL7jeChIWvYCqo4iT3PvnO01xM5z
UUy+vlGQtqv/pNh2EdpzyGdTxRiZ6t+Anpn+MBqBOQwVG0iVtMcWFM0CeKxULA4z
t+xeL4o5VUhsmLwdFad3LXAT8HHCguBLcV0/2yWijVleFZW3HB/rrL8ifhdK794l
EAEZm6zloJyQCln8K1oi6cm/g8jTzT1NjPB1N5Baujl9yl03ouyIPu2F3IFsBGBz
lPwo1HqCyESvSx/yU+HpiySxC7XpwYqP4rUSYP9v0uBrHbIXpHYF4baNzZ4CE0OP
ezGDufSR/moVdbtvWsvu+0CPjQFnrLLHTzfj3hovA5t4gsEKhLrg6M5P2bqw1RV8
CU0BxQGH86J17Xl/FCYjgkmRIeZULvkQ5Ajz2kgYrNxAsLfnqFWfPDti+6r95aA0
nzIy4SrXBJH+22YCovZcja1e8jSXPr1Gn1bGA6HZkJr/26WNNV0qPV4Rtu9n6cp8
R1pXtf6k3+pD0Y20dmaQCegtdQjo1OZFVNb90n5XgfVaHf/oRfQsYYciELtpTGpj
P5G8yqC/PVC9hhjXsnWj+Zi32teRp2jQwUbxi5UWBY4qzxDOPN5cg5qBOiM1b4zk
GrLJ6d+bkPYIKlsHLGQu6XzGvGipQtM2J5UAhkBHN0LWkhTO/RBqC0ULurvP3XCL
cc8o0jv+lDV4Z6VC5Q2mZC8NVGaaIVKN1jl2VWoJN0gtYYqNp8/XjDFjAACe8ZVV
z+aiIWDLv3J03ayU01t7u1ktiw/VBTITLQ/igoNFY7PFbwj2GCe3M8dZiWOUjYKw
ZsxnK0qHbObwENj4EkIED13reQ3fhJogz2N8oUMXJyI4ND30V1Biyugw+j8lEdUc
nl8hluSUDSYKy9tiwM1Gm8/KuoIJ0Evm4hUHRvfQ2z0ZfkNN7ujv+uFW/H27FnxW
JpoWu5a91FxIebE5iIhqSrlWaJUqQgezGONQ6xIajhCcOO4k/ZwMZN8hAHzFQ/ju
NimLEmB5r9LgtBQ9tCW8VF9l8qdHEVuShCkyoKWs5Q/8Q6vSb166rEOea6UbUFaV
9OdzMgn9V4jpVwI3e7MD7/OtyfQSbQOPMgooAGJGinOUM/NK9J82OpceQcdOB0Cy
diRLaESe8v9HbnXSiJGeYsDmNd7YTupugozH/lftKaMR6+kVEUEO6/lOxcyj0nYL
U6WeiRYvMAYT2mpjvv3Nrf+CX9d120J40YqB3iw20pNvLhRDoaGKQrWTM8JqS2gN
ioos6A+42cpICyJfJBejp1p6SxS1DocOQjuO9Lj0gOd/0g9Bjr4b1oPbGYccwZvk
/Z/cMXecBZU7mxDhrIUrVNjdHPR5D9WZ+47w0PvzIEIvxVr9jDw9HZzvMs5mft5N
8MyeBaU2uZMAtRlubM+/7ENr5jSpxrJXVdVUXlFCL3bpYxalu2uQKwkSU2n0yd9H
DPaUCke8s/kVsn0Eo0zPCWFIoMq7S1jXXyE5wtvj07VNMbrgaMEl6dKPg0S8dKeH
8VKQpx3SJBnP43/GEK0CYTU/PRqdAY6NurTN8O+E2v0HkLS3Md+wXx27Edx9idPA
oPUKaYBF2PUtR6TjKx38jOUbiI57Z5CSBEyIJwBsGpBIwWEBPyQsOAoSNXVxAvWo
VgoKAmRbLi9grBkzHnTVlNrrQGXHqJvf5UTwIDWzwGmCR9Kil6BvYiR2eOyyGpRH
6GlQeVBtWof0BCkMi6C/TFOZ+iSSlXs02H3W3ynS1zdqxIsR0YYpev0hBN1e+bnn
rGuvSbwaef3tt1VOVH5/TIiBJv9n2eN0V56cc0/GbwmfiQ8A1p0M56b22LmLMpnZ
Yua+NbDH+fF4pkCTQBabOKgiwAVR/x3mUk1soW6Q+Y+5/sQpCeyh8g9YZWba/oBa
RCIuP5xX5PUIascqei6E2HFSz81vCn59w7T562ki5hnfpKUM9lCdfTPseuGPkBNA
t18tMTE56ZCRnPzKoh4RpXnilsFwU/FmSq/my+9bIDqhB+9Mpn0lUVTbwxui0VHL
Uq7e7nXtD1nEChe/nKxkJsQeNu5vyIb80Peswq3O+ozcWd8OFba5ojtFkpdxmT7X
WsceULW2U6dIJOo/34IduvtmA9d0PPvdHhA0s7EXgqeYPR5Ap7CU/QVaewUeLaTM
oCRm/llLJftlQ2jQ3goU9A+M/7kIL/AJ6TSKs7jOl3zWnB+PJctIRmygaQpPQ4vB
lKMWg0bXoYC3SQjo0r7kP6nOFoqQPS7ucebp1v1MiZLqY58uT/EmOux5pZ5k8ka9
YKH1fH38Zo4hUirfbvwYIgJrBZv1q0YmiQJKpL0/xFnR8qYUxG3W3HBcyq4WWcDp
BfVVpFJ1aahbT6rRTebwnXZoeLY05bhv0u5Bix2HiFU66VtvYQVfv8Xt6hc2K8+v
PNKlEsMXgxLZsLw54qJXXEM7rDI/FDwS3gqrGHu/lWJaRCmcv9ROFp0VoS+wd5l1
PmINdyIYDCWkvCOEMaFVIp3ASD+SpG14c/WVjN0dkEpWgHrqELsUUKsyS6yFX/og
VfClAo5RSeZZXk5DAcv/K0ip21tSlukDIKY3fZB+k3gqS9kbc56UNpvK6xRej6gt
rse/2LFzWYEBYxlSe536oFhU4UPFP6m/Yv18fFJ3ayBLb48THVdUEchPmER9yBQk
81CSGBZgBwBa3fFRKK08SZJQZ3LZuO0o7VIqEdgP9rJkGJJIjM4wo0medGNdECGo
P2kdJ0pZ9Uzk6S2j661wkC9Fyr/hN5O9tfiT+LkyhvPnv1rWK0N7ros+RzkQXYNU
vEsbvFaGFRaL7NV6LKLm8gFEWutGY+1ViV0Smgpes5EKQGlw91lLv8Ke62ZU7Le1
mErCkJneSQvvDgvOzAQ8Sl376iwvTlY18Gz9vMstwZh9XQLUJ56ilUmItc3Bg8f7
wcgPsaK4x1pzvPA6kgzp/DwVe60h9T+Q+lsLvEMkw4vyufTSTFjwQu2Xtqr9k6AY
Rpe4ip1I95lV6rOBNo3tMVfXqTg0MQCUrI2hVaxjVOW2mVNWp35PSRY/QHKEiy+p
6UuROzEqR6nSDctsrceHxvUU/AOHdAOqZjYn+K7Hn1hU+yH4ic10HgQupH2mblSy
s96+RsKB2J7DB2fmkjtCPUIlcPeU8CmdF0E6PHO2I8czLjhaOZuQ2u/D9tTV/6ek
F8mTXwTZcET+UMHIO6XAxqro4C18ciqfKVMoWAUlg4NY1N7xhr1GX5QJQmahKqMf
wUPmt3MOlvENiBIAQMsjqULXWbMweeBEug2e0cY0FZXFN9UylGygST4soybXQHCT
8O7QVOzIBgKXUs6qll8pVoiOtSCqTshqL6n20G6VO2imRmMxV+CiftJ/sZwV+l3j
NI7Hh54WNyBZlRghtmhqi8CWu2YSL9FVDJQFEmFIXyQrWJticn+KZFdP4lpb1Os3
1N2MW+HHvr1coiSIqCxDqzQ9TdGCgChTpDLw2SoVEJoKVhNWWS5qxq+jgAz5p1wj
XgOiCqlSZSa2xOUXrDOVoyMiIio5j2dTqzEQQeuXdk2SGDFOvwVXciRbGIw6ymDN
9bGZ6TtrOdiN/lrYXMoFlhi3YbW619lY+L0dtnnjbRrNkXZ0kJxDdbFY0wCXvDhF
w7V+mYJrvNnJ8QQny+Qmor1GYpW1xSt5KTxpyvbpIpmzT7TCfN8JCgp6Y5mW69WW
B+CrdP/ziBmbvWCoNOJzyZFlhR+Iq54ItttKcVQRoQ/OJ4OjJ82a7PhXHYThGAiQ
TYiSgZrdTd6MuYDssajmV5VJ0Xb3MHkWLee4Us92cW+3zrLXzqP3lQ961KGpeMTg
/7i75wbkyNzVbaF/UNkayeiGiU36hwC4eldk4WxVq5w6tm36D0kSLOjf7N4Pf5xR
NZij3wirbf+ZWonPdUL+iQ57Bw6oQzqGnRh0WmGgeYuViHLGLCO0h1QD8whTFoq3
LxJ4QUyGpb6miApeNJxQL1IC0hl+qkMf4VK6GpQAIaYJUABc8JAhAAlJDjYaoKpx
5jCmWhq16M5GFkwCDkIXq3Px3KpVbPmRsXqrA1X8F6tWtXsVsFm4WGfgu6aWi+El
TfwAfzVHoeYpzuYVXchBtbjVtnGTaC/E3q7wWs80dLegTMsbW9BSYLijMlh4L1Dd
RrypNez1YsM8szdD5HAPtA4f0IeBzgaIr0P/G8LnFZXGJ7CSwxAP8xEVoma2fL0Q
B3ZxPLgDYjdRlCseOe6CJUk2kGq1Z6YefTIEUw3XO+IiC2VgmBveKHtKqjFXJXfy
STp/HyTGz1IlYbFwpnXFEy4nF5qxppIlU4ENBTVkqE2whPxXu4Ig8vzOYLvVVDgK
4hfRJrvNm7FlPZNO6lLn9IhgbXik9twUKWL7+3CLB1jWxRAfskHUjcnmCQtcOXDJ
uoPs4bslGt6dQALApT7MNS/YL4gBuuRN7rQ4YHbnC9axa4H+SXt5xFrGRGJ7uCJX
3kd0QcOvt/gCi3b5EN47fTM1yBKQYZA+YsdIvPSiBiVOW2ZQTZN2Mwu/F1iWgqRg
jMu99hNufFAH7mlrkvajy2RIQEXADSgtc5CdUNZfM+CBze5shLzW4wiVxV+uXOGF
/6/KiOxhokU8LGh+89+FYiIQNGkuGPIlklzGThl3gdzcoKfHO5kKv09NH6UnFcV7
DJFKtjuHsqMvUjnQaVvqRD+1YOhnthgZxtz1IyYsuQ4fyBoGmrZ5MzKpixQWm5RV
9lLp5ULBiv4m7USyjO21LHwpiwLbKR+juIMzgwRfkZyCjqB9ufIZVLDop71ALbYx
I6aVHKq577+ybsrChUmIXa8pJjnHZey7dnT+3GGaxLV6yQQCW946056odocBWt7A
b2Ob+4erYhKMkLTazkRx2cHvZENHTjZETIJocHV8FNHWZ/g2g7fx5KgwknFNQB6b
/4or2MbIt4mYCaNJjdgFXJUL6eI+6ZjDUmPABgGPOOUJfkxkuor7zM/VXSnnFKBV
oXpIGhm8oSxBGpSvJzkhWQAClPRCb+CyKpS3Q/z/ak78JecngC/JqQr1c9jjzLlU
TTKDfZc9OI3BEvEGj5q/M8ZDcQUwYupon7b31evAU82OupHnLlMOckRcuFCptwa1
rK3SY/TWvM0fXjPxTp87EU1m4ZDoblmo++ev/ADYwUiRJHPRFvCS4mBFusV2xoAY
tmEeXrmpYOSQrpialbjscusBYXx1+Ev4w8hEf7t8AdPpVAzwXdeSoSoiD6+hnhpX
TiNYPapK1xwSGrGuWBJqtU45MmFTNHm4PKMVLkw9V3hQzgkB/08YhIF88X/OKYEf
75xFtVcBrflzK6m7l2sceFvdjJezljnA7yXOLFX3PJbzuTNDgjDzH0tM5t01ypQU
if7JnIWp11Hbls6KWJxVLwI4s0xWr+MGNgtSTdJ2pYzSMg7fdJeG/zfGx4nhbTEF
KCuEm2KxqiFkx4rJl5lRNOk1XRQp2rfon0n83NNSDp0ftW0UMVkBBB/n/Z/OQeAm
p1PlT7IJBSqlIReFthJHu3gtuz9nufsEpbc3BlTWRzAELzNH7jNkB06PmizU1aTG
JFVKk9GeBKdTZI2+l8i2XIBjtB8nUIV0FBrL3AztY/rcUoa7JLapLAbZt5/kb3jF
khq/3z9SveQCpLsJc5Eq7JA1NGLeoUteflyg8MHXhyijDs2t8pq/XlJSujYMhmSd
3EFxO3otkV5Oypy+hEg+xlnS1TbGPb0KvFmylsShChwvGxv3Y3KE9apSQoC3wXSJ
C1Q+dPJy0kWDnolYy+HVU5YEizXkeIc3LwKy4c7VJqPFXqF2IGq25fmiN80y/dRN
iJC8eZCD/YJkpuiM8Uj321EwdgKWFcBGQOku79sclMu9WZ2O1jRZmjGvV2gXSQEB
u9rfumUeraEm7T1gcwPVzbMNY5RA0I12CRerJG8ExXz+c5b/+mZWSrhnVs6uBzHE
TtgUDj1jq1uYDe8QjhuaRQh/4j4KKNEQydQBRmENbmv15F/vVv30S2NLEJz/0etN
YGnuHObTo99S/Y2BR9gPmokL1a1DWHMXngSdEkBb+SLREfgxPP3huZHRhOvzApBZ
c2+RV3e4PdigxDzOI/i11MY65X+4EmGmvW62Pzmls+gSUdMVnYeiSTFlLqvtJP9K
eOZpMkXBY8kzd/L9WFN91VUBxA1pCyqZKgk0QJ9CfDFgI7TqM+Txt81aR7X91Nt1
CIhqY9fmyPxMWC7yyAstR1aoud2wYDrV2fOyF6/GPpbwaZLUdzeege9xctTPwCv1
4V8xPObaAKSOegkHEFnS9aLFzr9FOfUKZO06JKhSR7pkLTJTUPwttkbzV0dD/Was
m3TQoNbL2YZ3XS/tNM8/8cv3e+cnvZ7t+vL4LrUAfB8q8bTtWXhRvU7w0dc4QU5p
7t65Je4OvHAKKSC5vzxyBnT2ACnaLQHeBResio2u71PzNDnEcRtu1VxtqeNFJNIy
Wb5znB12FqH+/aMcWMJRMLDh0r7KuA/sy3zNHsYPytd6IySQcuJjY/QPg3VCMPZq
vWqTOdjrNhTzT6H4Fc1kajKi/Oa5CUpQxKoEPrB/NBqQ+BK1t537eVSz4JBgsHEJ
qtRYT24nOcBmAINfb4Yar2n0YJTUuMBoHJ4Yv4dzNUFRBbjKNGeaDIYL/8ZDECmJ
osZNcnvOhEpkhupB48FPLmvqg3Y//gVWrE1wVt2mVNpNgzSjRcR2/Q4D65CqB+Re
bfaEnmcrBBkgcK9lfGWTwTFlsgqCyK3SXE+uOyTTfah5XcceKzTPX0tbb7fAaLap
SMOLcluO0zLX9lB0G1r/Ljx/0JJV3+hKfPBRjBILDQppMT+WrTAOHENH9qaZCKMS
i0Qndh2GYBSFROiz5urVADqpbky7lQ3et2kT9rgpCI3MU0ghoHPkY26enE0mI1uf
EIU2dnzin7H9hZwY9vPzWZb2zSu8yqU3I843l1P6Tox5WUta4FOvgVizWyPRiO2t
RJ5j++FSAvQyH3gCQjxw/g011+e/CcB+HsYd3IU5yNVdtpQmvKBnieHwjLeVWgyp
zXPLCOhRwAYq6IMBB1Yxxk64AXEia0kfo06bfv0UcFQR6jv1Wq3sJJiCpZqYhTmO
lMJVKaFeRz2POa23fdx0iCQAt4IlEnR7VyZ3Erm6IwdIhrhyVICik3DNyXyiZuBP
nSJRWy/XvW0N3I2FDiaHCD9qdE13M0cXrbBN4LPKZX1aNXAcNQTx0NXU7OJ/Wj1h
3rbz2uZ9D2p6h5HVVMs7ufhe8ionXcZGeyU2IVgPMGR8IwRQa9GcccZnbE2z9KkX
IXUccbr+6m5P30jDHeU5hzah/T5Mija784iZ2B1uBB2na6HdeFn0hNXoCGa7RRI6
mUkru7/osSUyqtGfb+DSlLZJyLlbADOpfSNmhS4bEMXYpHXOlKTWc05AN7VieNnI
PMU3rGHXqKr3KDwhair2RgyKm9IY0El0OFn04rI5ZmS70QLVwi1zn8Qh3ZbI5Nlx
XxeNkqBCpK/qZhLb6+h65XHg/ZIWBdt5RmLNYjT8DQRwj++bAqdhwftmuAUZg8rY
H0EZN4AVRxuFZko4PvQiiy+VVsbk5ZIA7CNwVvIxn1WJ86zyWs7e3Zp15BpXU6g8
t9JDqpcrierwnk+0ybVrchtfHbYRg8d3mFnCBpM9Y/WShzCIr4OP6jdtB9eORlkf
ROl5z+xHnaY7dIH25ZbjbvrQ8nsqJczMQRzr7+vBFZLqwxlB9HqoPzqL7ydx9e1D
mTYeHuD0+Qh/YbTZmyFnh/TSize0UI3bDouj12BBA3QAQ65aL5mkAj6eRSa6pFU6
vc5z5j6RlqQJ1nedRv9jeCIEghaJM2A6U+qFac1zyBLs5nleF9sL3iC2BJqzLgVV
o/OcoR6gq+ZUipcoaLWXOaY0bhHsffETpQVUJ/J5EgN7TATXjScz8JLswD+4QaRH
YVl2oCY4LcPsUJaFe9Mov9J6oiAQqSH4p0+ULUWdNqoVMzHOeRzwEVQKqCbpWs8D
qMlTk0FMsIcIrE1bH5wps4szRBGFSXlQp8EfQuHYtn+2Rts6dSGJbJ83doPjeV19
722pqo7wbgCOAbs8QJ/Ia8IzQ+vlDLg3jGw8jk6pkg0hz/c5r/tZhTkP6UOjdUiT
pbto36RJAld6DINUPA8ucaSM/6siOCGDHDzdAJ33EsbegJEE0fLEhU/UyoeuGSrA
yn1V5+mVHoGgXY8IyLuw3FwAbs81X8vqAwG84JGnLEn3o0bTt4t+elmXxJnkEoG9
OTuD8cpMgmhY8rYjGrZNee6lss8TkGcEWFcL7qUt42f/g8rjTm0/SOgOg724trvY
NEbttyaYjuqpmky2NLy63pKZekmXkIxyDN589kc/NWk/HkqOlDi9udHc332KNq50
Kc64D3PROd+0E3YbD/W7TWBPLOrtm76ls7eT7pHtGL4uT0WSfVbe9PuNXTHQZOwT
B1G8iXVhmciJ+EN0/WN4kivB6ChDLnMqUL2tvhbgJHqe57KsC4yNDUsuwfbfhY2E
fwmUGx2wp45x5CUaiirEvZ61Iw3OCeFmCfCnczlJYdazUjy1RoJlfeWyBDqz0DyD
uy/U5k/nKdQp43jCn9gzE7UGpaibscVZEny/MG8Vv6N12hhaBfm23ActPpw2UW3u
ePdMG39ApfDBItbJ0i0t5GBlAskQcw/kyVfT5j/aT949gnrovhltdY9pGfgm3siO
QqtjaKumXB18U8aBxOQYkUYTdaNshhLGnEVgtwgYZTQsKpP3MWlQcE4N13xEkdYq
lKuGVknxEfSHYWUXfqlteueHPdVRBZ2X0IHtO7dJMlhS29ZJpduD4HN9lTE2ONAI
iguiizorWHKtqCQiBIi81U81oIo6EFN5lMRGt2HrRnhtGezlf+cITxbhnDeTJNs3
DeJp+HTH5qmEZhZszyGybx9eZIT6s/WVLi0aqgG0Onz0dLkN2HOj18LPG8DOotOx
J7PKHXH0pZNBCtnEY237YAB1FQ+He/w+67GyYpfzy4ItuD7P2Nd2v9/AOPA6RfVQ
xwN/ggEAJFf9rLNbDTLOMnIXxfaOEdfnE7eoJV1dL0fga1QO6GJT59oFDkd3A5jn
gLzi6m79hNE7Hl/xA3q67CChUCsIs8bFB/cvRrgOhx2DPGSfoXeSWoSz2f0vRH+H
+Cqtv631OMZ5sLdqj2SK/XjebFgTTLX5udOu7lluW7hdqhoGNPufmkVT41CGl9Y5
7umPAt/k8P8wUZ4owdQvWKYGZzTSKav+Pjd7ixFRqbvwZen6qeLVTRzztJ70DpK1
QVXDy8Jc3kQWVNiadfnpCP5u9GzQHvEJunT1fOau8KKrlT5czuaVA+ZXmO+LVA2U
niIjJzgnbHbX87NwAqWTAIVNFf/qBAM7N0puBdbPGLujU6TYHmWkbHur2YpswGdQ
R2I+eAN0FMA+5RtNGm9qhC3N9l3gmoCh7VmSFQghEaBzzZrc86kZSEwocaZJt0bZ
E5R5yKWhynNEmTpwnz/DEyCQZh52Ku5cszrMGHrrFEPBEdcQDFQUfui+XOJUaLYU
KvKMy1nBtLKEYJZHIAe4zpNW8lcl1EKRVTrC+VMJWhzE3j3ra7ZVW+ighmP52bTj
ZtHZDsbwgto4CX/lQuN9tZ7jYlp0Ne+gRec7Urk9tcty0iO7y5wDsC3PjH3X/3OM
GFT/RzREPr0DXnarsRWBEHYzuivw9MxgiTpXfyJJPiQEXInYhkWBTuPBSdSRDi5q
87qmvbkkcpXn5qEx7yr+oTnSePl/FV4RWLnSq2kekv79QhblG8e2akxqLvRdEI6m
+kd4AjGuQjAVQ41589OwGvKijnlT2nxntx5Z7lwWLenTJomwNmi0eF+O1CZ8UwKs
Q/yJThetztQnHl0LdWDhyugIoC/ZcyOB3FWoax7+zmYhBCtYGHHfp/gQZWNhxEt5
e7CZN3EgtJJAYCmuKh0j0O80usdk/SEZoDHRQuXS8o/xI6EoEEiOQo3n2z9cl9qX
Evvz9duPDNRj9Ztyv+cuQ/bGMO7DZAi9eeNS7lUjfDVe4DtRxNNnD1SHiBRzsYW7
HzOVeSTW8GcfGIrOC+JSRWixnlN8UreVieCtHiUshSXKAMBeC0Zmx2lSuxdqtuta
2ZAem63Kz1FcSC0q+PWM+28clvWiAK9A3HuUxDtLPx32Ou1RSh+2thtMYh8LLKhM
+10eEsHDz5u2W71tv1SFq6hoXUDJupfHIc1w7vOGUcDMoem0dFH7xwV1+xqCq8uc
5uECU0cQglkzt1VC9SHIpG3HGZXuVnEoa5JOOFQapZGW2liC/4SfS4n/kUSz3Xkw
LoFxuqUhF6B89kJbC5dJdzavN2R0dqOoT3pnkUCrddDSSJfIcRuLyWf0lxUWkSXg
ndmftFAPfnzJSdtvB8qljO5t+8yhWlHcKMTltjDCnWqJRuVj553E9AB5RO6hny3+
d7KJrhvBRAQppGVQSEmhN3dvmjIyL49YkJnhherONxpjaxP+Waf1BJqpWxwB3qzD
lbkZFxeItDgNkRUJg/VGPct/iDuF2V4Na8FKi1/j+8O816dXEdELGGz843vWPfY0
hFBd5o6hgCYl+5OzSe6LU3JYHj1KIbfv4Rxv3Sx3s3+xEZlTk53c8SYjk1ce6bq4
b7VkDlqqb1h1bNeAj1yj6S5pq/nTDMqKj1ksLtf00BAiL9EAwDeSaG+GbFjPBrmO
ciMlwkqY+oXyRmVT/W5AOggq7ligO6MgIZCwCK9NUBuvRAudJYVTxVDtT18BSz7q
3tLxgPh2QSM4eOEEbvZ46Kk4Xh+e1Y6OZz20QLSc0aw72O4QogIXoElEuO5Uvso2
ZN4FczMdhnirlr2pQqPjZIOp48G+iMp8Kg8CwE2k4hhnhxbTf+WpG7TRgPF2ns9i
jrK/nxG3m8kkwQHLnQt0CYlPay3zPpyFhTGxs3hcRJ8u+Xf5q7BWEqIA02+IAqtj
taj2AT0WurqPkcx+rLjIU4v5UNzcTLL5vdBZbPMyY+1ccfzxwz64lFokb/6ehVAN
Zf9+hsugNYO09UNCDprIciURdOISxeOYVqF400xtzV3TOffQNNKCLiOfkxKYsqFd
TWceZaIQm7QECcDH8rLpks9w+NNQIvC4qMs1z313CH9dNn8E1S70jCX5jVwJUd0I
SQ17CqJgGihlJpsLY+LUMpbujzJuclevZj7DDXRmBbueI0P0RXny6vVkzCRM2zPu
VMbhq4JjvdAlbHltxXWFMNFCNaUOjfPQ/g3B1Jy4WIZ7pSaSEAsvnZacDVYA9w8T
YtJrgrTxA6h/6fEHry7ahGfIWr0cVt6ROiZ/iScASxwksrQm1Cw+1FL+dpFfatui
sRwGIkn12qOGeoZK0uUwsn9opRQ9Xpk5Awpl8I2CS9CCWiBCqyICGaghK+NU389z
qSvsMcviW9N4KBEW3nxb3xG4PUK8w6KLtt8otM+W1ScY7S6hAhFodZ6K/a3uQLQ9
pLApMckrpOmBdjokF0jolMXF029AJ1gr4rsfv1jO9G+UlULFnIfYB341ISceLeIs
+kkdPxp/g23m3meYUxjaUnralZ9A87irEmcytTbEa4GnZGgWIk8ecPVT49asZcsB
ZtXBuMmCgoHQMIEJ+WlLz8HSa01n5zrHSYaMlsQOUp715Oasjsjuruut9Y90WoYY
T1uujKauhyfVb1tACoODX3NQNBZaW2z1mIMZUhLuS6HuNFRpB4wJy8GW4gjORcws
2P5Yn+ht1Slx9DhoGBb9BDUoy2XjzSoFncB1n4pm9AI+RXZyYd6akb/V403WsBNm
AzfcM+FmxZt4EGbUETRyP/sBw7SpL9Ubez0zhcawHAlQensTJw7Q+EAplLhmSBJf
L1umbd0hTD3sJeQs+Ery0hBBdIIehble+KUo9DmIQezFWo07EsQwBmtSFeXBFkiT
qKnyanpV41KFBG3oHKXiKBeW7PLH2Rol9FD0hIHRwLThQ1blXTvwRpTcGu2ZwUtt
kQCtmkr+dj2WMChJa7ru+opPu10Zx7FzBNVxmnCnsmQQDmWAOQA2TTYol5lsqEsj
TauRnIAte1cHKGMeyjzgSeEbX/djPb/9OqWCoUkMYjuVFcR8D6PF+32HKgrvUQ/5
XhKR/cLu8pUBUQt38DKH4kFPxMI0lZRZSNNd7pDJWHfaMub/VaLzmuThs+B1nmsb
yqffU5DnTdymRRg7G0CXiqnAB3hm09nECHmgpi/oZ1ye85pYjMoO8t7qyTbEj7gd
9F75I9WBq9Twz/WfWZosXlavvRsO7ZRfmzMQz7ysmROxelt3IugMTA74viRr9Kun
I3dn7Evfx9UsXXdXSx8hDKITACyzwv8Q+hgWQUCi0P6bqhCT+zHIyE/nnDg+vaWj
8ifVV3Mzz1R0lAK7LxqG4Cuslj+lQhDJKzeGh8cW3JITw0a3WNx3iH7OUhXSAvC0
1JI1LVKXjFK5UIvL2DmJ3/926DacQWGQed/b/v+tF/SQ1Koq4GPo6olgzconiGXD
nMjXv59+XSrGJ2xkCKswUw6QXBXSpBxDBd3XKUboobj2xclDcYuk0klBBN+OyK0m
+PWpMe67kwCPP7bche7yWRhiz5s2yaNaYdOFHL2BdrTLvmLp9bC5mVY0zDPrsYDD
53FF9XTC+CFKQ5+JxWvaOHGhDEMcOA0lqfR7qlw71lIqP05KiFiXynGkVPzhYOkp
6p1IYrK3R4XR2Id4ZF9z4DS387POnZykvgFmHgRIePIqL0VVFM4EuuMM14KaebfU
PiFITSVLWXJy87ITygi5ABzU5nGKzU3b4jWLaog1NpwV4o2/ZYzUXZsApmagcGyO
jBVZyMc9v6ostZdsGo8oZNcgfx1es/11ouXBzK8X3oE0rQvhJamWe4MbBI34ie43
5r706mS06DJH6owjiQjeuWOCtVi0QQx60M7WwFZyejSSvAg0tKzHOMmqBbebIInt
3kCvw6/Xy8fDsTHdN9WENHX9/fB9BBvw6G1wH6p7ke//ZR1AIjQuFGwfNRT6MvQa
bvMvwKlPtmopkR87pSYd9DBhKWDOGp3FAJxYdd/hgXcOOV//7YMnzovLqlOuI1dz
QSqX3q89JwTIX9mYaxvQKHLSuNPunpHYaI1biBs/gi9vvKaCp5/w8WpzmarO/hv6
juvlBn5X3BCK6tMlRkMEm71uT+Cw9uoam8JHwjk0XwT1QWaUSHqXfeMQ54nCdAU+
5rOFsXfXBdocohr6rCakI9smIL6W7lCZTscRjQ6527ZiQJn8ASy8NNtZ7BYVQLCU
CL/MHC60wkiMoMobLNxHCpwciY3f25F5QVoRcOd9i1ZG16hko+pSMb7h/8DTGk/+
ZJxePBaV6TZjODbDOqcpFbs5LMzYQkiLEU6PmOecu1HZlrUx1vRYkVdoFLGmj5xR
DXHFXrg4boO8iyQbO/8pVDWlDnMNVwYEpuA+nkBncQW0uDqONCuH9PXidt0WgHdm
PxkSC6Mq4dffdnPetzc/KgVcoao7+3t8TTahPkjCFcJsOrIDPuHnkcO2NB0OdhGT
iDPgBNTdeCVghdY6YI9Lyf4nEIj54875ALArTC6yjDBvLxtn2U9CXM6sG6B+GNbl
9/qEAI9tM2ggq1jKsBObsDGV73WbvhzfeaThQtKLGcPA24M01w7j5luS9ImLEtQ3
tbA0WbNp5pwvOEdgxlPeiTlnlZw/ssuMiU1nwloa4wpwtUbGs+Ja7dVi51FolSTB
WaZoeUSwJzgGUA0iUEePusF72Ba2ztIHNXLZrjJNoM4vf5KTEkxF5kU801crIYFJ
Qfkt53S3mNVwAkJ1ZbalwGVo7eSHjh8B/09V7+HhDwUcmICv95z8Ux1YHT9rIXQR
oai+wVGGkyumfZEZ/gaNmr2A84jU7zxmXDk6kmiXJsEgWXFF0+aHOjjgCYpkbEeJ
W1KO8E+Qx/v/R9UkssDihTh0F889qlB3vIoHRzCmvLHlVkxgN9Hv+2p1Pf+VH9kj
ssErTnP3/PWfn5L/AB872Ir9lZW3d8wj428tRiNVhyOC+M32sdnU12ghaNV0FSlc
n37lmiZ1kSzxJPNkD+pN/uF6XjHPsUsaWPyQn9G+0huG2gBavUF4OAMKFnuNzBx9
PTBwCbcNz7AmZ143nsW1X7qq7S8xHfXUgPRD9VLWY0dHRO++zXUhUTj69KOG4UH0
cagGluRpipkDOrFvDISWW+2vycU9pMiTJxTTHyL1tJcXvjIUbqusM7Azuq7qHoz6
h2/QfL+cW3hMLuDq2JAbrkb3IlEb2aiM4Gg3nXZ6Rp4IPt9K9P06XFEt/0bGB4aa
hX4aUKpz/1eRlH6Jl4y3kgjHibneadUhC8Su2XkoUS/oCGtPaODAVi1XVu3hwoKM
mYJg4/SBi4KDmk9AJ9wJ34Z+/pFxVRi05pqkFo5dFsf7Arb1FSw2Rjw4nIt5Xek4
K/VqxlvoxygKGWLYXXFEDknqPfchee7Gn86hZW2AtPp+wFjb7tteIA8E+mxxEMmW
pgjFms55lfIaDlA0bl2BQB/AOjqzzAtFaZT3xcw+R3zF+gdiq28c1q/DqpL4qNNP
lKR0xuV3i6vsDYaOG7MN6wcWDZ7KS6CJ4qXsSF6QtH9pVTwRL+KESkP8QNdrZj+z
Fk2Z53JfiJGcJe96TKm+jyoHxZ3yYPIjXW8OOuF6eA8QayVsNl2vuFMj3Au5Ti5G
pD71g2j43+3qmVpeVfe2I6xj9ZgKgWD6W5UnaaWVeggzoZVu0/fdssH4qCm7Pqqt
+bQ80i8iChZSUHhGfWIk2HqASZrzQo4xdZWNjMQEKbSuuynQ1wN1dbi1LCa6NIjQ
92oDAH/W9psr7hCHlDR5s28ukuGHblL/MnDZ1cCRYOqNY9ZrehTOMomwVw45I3Jj
0vroPeTBd6WCFRLCH1ZOHmtC4lza4yUy3oSho5Fa5gHzWVM/9S9JvTTKYQCcmGbs
jwjCddr1XVA2zzdqkEjp2NusMMS2gTspVh+7p5per8loORtpxmaH3RCK462DBHtZ
yXOFlTrHLhzi/jwTo2h4Gs4zl595vb9pplOOJoawEAlQP8wYf4LN627UsRjl5kgh
u0x/qQATAblaNanndR1qxbijEh1IQB6RazbWGJTrbL62e+U7iPaSuhQaI5+gDNgc
Fv2EM0MMj5Kek15YuZI8Xt4UcK+oVaNnm4YdYCcTZAkAO8COvXnd8+U40bjDK7Gz
6KHuRxUMsRC3rYjmB0ZxHkF8t1r3mnE1oZI4E7KkeDV0UMGAo8tpocicROvf2+p0
P2ExU6t/MVq6Tvf7USw9Lbpz5LS2rktO9u4Le4ezxeJFig2t9ZPWPXpq8bIR9wUh
X5YfiwJAWXDQbb8/KxPgJSvUoz9rjWhb1g3fMpxa39WyKLa0Ueyl712tif8VfhGO
hCHkzrCa3cmC4OyeYQtRaFa1A4451IwesxtOXwIyfpT46eZav/zvMwc0jbtiB5zu
ZXJg+Rdk15twHxTLh+vYBxTnUl66Q3AUbBTcsuiYLot3uMWi0RKOG6Uo+E3BZccS
+mojuwDUfqlTKn7DblueEzOv/Kk/XY9azg3MtqrQ5wOzIIrqOcrLoBlC6cUGiByn
zvFCdURuOZ0B6h5u+tgJMI8RhIZsD09hj28TCL8Nea6Joj3poFfD6mhGt7E+aLa7
DrucZFDzBAKCg1/y3nWgkmKcL7OBxu43UAMAqkGwaXKex9kqi5MErJbA/Ix7nXJn
zSaVNte+R2gOwjLAWpiNsglKy+MSR7IQvjUZVhqdamD06jxSghlt9cCivxyJmZt3
STzhnZul9jDwgdE6BWJ0+9evVHf7WxbGXNTCb927CVWdIgxwe4E+MQVKanIwPThE
eYypCnRkaLVFimK4vdf1so1hAUchB9yFnVO09RwbV43FpZRfOhPhxbj2dY3WuDr5
Z2kNrVMNP3IcCMIPFl6HM2iBvUpq5DB09VeTGtI5kMyNVuAjYzixzEG2neE7OTr8
GHBLG6DjHq06lUffhAOPN6m3PLdJgW1K7wRK/DWM6nRCeBvtRkw1aOolePxQhF0G
DYQGpzvTrfvZnDLivC610W0T/XJAfycDEVzVk88NkGGv2of09B8bsUmcsHl4dKYz
ZysZzdo7E21En/UfQzx0pVoUUlBa5xFqgZQRyNRJADvoXCUI6wuVtYnOeT1E7Bga
dG/5bKGBEvrEHQ01eeG56advsrbC4ZEtvIyqvNDGcfkV0hrwt3EpJPpZAqJ3rLtW
wIimiJ7TGGtnciDPPzctgM/7M8XK1mu8CRhDW7V9ox5D+EFjMBqoOzTNysgihpg2
0SqHQePeSlXsuoMVgffujxq3aRIpUTZtSG/mI8iZgLCLSArnmTNLp5derFtMUZ0c
ZYQ0W7lAaY3MEfKrml7XzrNQsgFcinDfe12JoK6Bq6xQ9kHjo4ocMqQT3YeMs1jr
xA5hSrYW3QYX7p+mcbq7rdV2JSVsap102lWpsz64p60qdGJSHaSCjz4wGHT3xztf
Q1Qi091WXfT8zjr7tdPYLfCe7eKP+RomCw10wmvir+DCIf51TFaCqbGy3nZdArA7
8bKlXjXxpAWKVc+3pOR75sPXfAX1ddzH7QHPqvSj0Z+jJowsbOpz9VB1d4joJaY7
4uF8Rr4dIY/v9WiJGXR1fjCruwBJQ/j+QM/5t7gmweBGmlfyU4jQgFjHEv4v0Kso
27NY65EIKwMhfN2xuClbayI2GgO1dWdeG9AEGGDZgKhbXNy5wmR3hlr8rd50iId0
8mZU0p4zbN+uOmIiFU+gtHHWluTFc51mpWE2iEFskbSqayxDaXepcWPmWw/yTS/L
dZ/G0ySIPZNvO8s3lx2oEe8EoZUSaPMW/ituOGz6+hSOwgOV2SpVRJdC5LE5AQV0
IqwI/XO6y6MbJK73BDtQdmE4/tsf1qYB1jY5Y7QgGdpiVQxhyaBCaf11RDzIHP7d
nKwS/GKCH//WAemIKFCQZr/4mmeX4OH44od4aLgcbkA5yxyAb7v7C5Gm67J9IY8V
RSs9eDeIFPEX4xquof47/iKDALI4mGz7GFXXBs6W67HHtHU+jBzOrPR/nNfpvKvu
eKmm1pV58y3HG/LFkFX5q0HVU+zX/RkF44XLRtwk3luSda4tqecB4DkIyWof3i0Z
lBkz4GqD8m7TInt9+x7eE5c3DXZO+JU99Pv4fi+o9hKwjsZCS1iOmYxauQ+BLF2v
gMLAtVSapHzt47VgSRlJZIe79XH5L1jZRroWfSyKOOIi2Xs1lm0Yxg7gzWshDw5Z
I47KnUwh8/wHcI+x+yEzq8pmtFG3LKd90sHSfjHvovUWgl9+7YkpV48YL+WoQhdA
8mC8vPFF0CWfHcYv61DelMUNg8s4S5xGMupNtOQRN6zAStFNf+19OuCNvjIdzq+U
igUaZx7TfNdABEXV/t5srYFNgBsJm6RgDj6uK5Wtio9BpQIn/qtl5uumYyfAtf5H
6Xhw/WihBqeWn85D25ZurVtHpPtRVjdxN8AvI5jBgfeVXooirqQZ7j/3o18mmwqF
FfautYFQNx68fRCr/+1cFQMbi8qWxDN5Gd449zEveoIidEIDT8e4FXh/JpHzstI0
xytqD7yy21juRqXyg2j5325zILH+AcY2GqcRK0JHkiJGkLeFk6ZrvLrfMOVn8ZfT
RrakRWqtvdkQNRguuKaMIGRWBIzwlE9CeGrn5MSfhP87D1/Sz5ldBvt124yHy47K
MND5sNUr6N0TIaPFCIel3AggQ0wIv4q/LBaw8phA6eGukeb3Gs0Kwwt5O5R0nOjV
XBM0OW18RIPN9qmA/vS9uU8kH2jK2Eq4g/ztdjv9SeM6rm3hJr5u5iWQxWdtBgpm
ctQg1GObv4jLDvL6pfJnEZI8ienpfiBr1BrifktWxWgEyFZBHn2EVyMRlDL2CJ1Y
ErGmAZUTwUYA79vbyVNRhukwCqUaWoWZapj1hx9jwTs4xGGWZQrHtvVjFlTm7CZe
E7xhL3yo2hxfa45RM0dJixwXaXB8yiOAyWhAwLPwgIKdai3wCWWhWBNP2ZLzqM93
Lq0XezgjoQW6cWd58OABLk4Dv6H0T2HYaC5rL++CVbcBAKZY7L0caeLnRDEyPKHf
nP6G7LmqUobQXijhzlMbCHXeWqw85Sqa3mf1aUo0kCYWRQt+JhaVCKfuN1vwVPY9
PfTyJyjC0hJlnZSWifJ19l8ZqixDZksL13yI5cfxObVngKum8U9LBb7Af35FDzIf
x9/AyOdVmloIDVPhlGEcdyXpmkXg9VytXM/FjWQYAWgMsP0cB9tGgscXlMMsIWzH
/IeQ13c3DpKHoGTKZs7Oxw1k8NcOLESuZwjB2cMmXwxL9jAm1UkhzAELZoO8fDdS
eZau8Hwxd/r49NfhflvVxHPZrr+162DzdbcOAyqbaSSek/T7kNSZwS+1S2xF+/zg
vb6hlXeifuUfJ8ubKiMVy6CuwWwdxxcYA8XeaWMSnzMYO9MlLp4Y0W7hN54KvdK6
hWEv8LhtID6Jw4dMymCAq/2xi6OPyewCMWUglj0wlxT321/+SzQoAJZ9zUg0mGqH
/BoQ6KwxOOd0eEOU8kHTNibAmHklaMr3CkYZ090rAe4XxPuFOr7lAWEAoqSIR406
PyGH0kTb+j1kENEFkrRLZV543UW9t4uSeRO+k4EL9VbY95OvsZMteu/fAC0Y/xOz
UdE0l5xBekb/oS3srIc6SXU3oF+nRVMXE6TGNGiL0Nvj4hEr6WYJUxLC6Mn3B20N
0z6RYnsbuCP+iiCL7MQmoZKkPqub9OWxOnOq0QmJ7WqjPiwZU+LoNu/kZ+kYEcsi
+ezuFG3X5ez+sQdoTxxF7BCqZpXXQupZnG4D9ZvFqAejEqWwZ0qNV4HWMen3R7u3
iT92iIE6lw0N1qKTFrsPpuDcn2la/u84l+KmyprOLJqC5sc5a/vnTQuYMbUbKhuD
rj3hH3ORpBbkvdKZ5bjkxO+6AglVDoWcG62HjSbhqYycve6mp1/nDmI0yPu8kCb/
2g7owOuIAjgj+imAE1pFi4Aosc6iSMXFgnzYvQ9L/8HTUR8KKYtbR7MuCNF48RYF
jqzBh/XAH9Kp16BvJo+DD5wvLVmo7bozWQEdnWSqcXwj2O1cnf/KJ+eXSwobrdll
cXCgF98STD6RvHY+PAUKhOVVXYtKg6pVWJWz0JD4MKyrDXc3OsKg21rHnfG+3Dc/
g6Wd4Xe4SDErj3HwxAahcqzHqrcYX9/cBOtiz/8kCm/+0gMBK06gLxTMS2W1xi0V
CdX5878oCSaJwoEggLFfQNCnMoAOSJ/15vDZT7aUQnuXM16iMbSU6pv1r07Belts
9I50eh5+mqtgIIWKGg+mJn6HpypvwRzOvoQyQ9lZSsK9/AL1czkFzBJ7Ydkfhw/Z
qxRnCdgmQ9Ar49rYaUcOuV56fCB6m6Kzq2c+AK1K+00pQySwIv6kBj4O35/1ruJ7
0El7CBj+uaWkRV3z1QKKjX5HxY7zWSJTjhbSjZ3/4CUNnweJe4X+hhlOyyW+aK9h
qgzRBO/wMqN8dwNfv1t/0ily35lmeBw9PlFKk610GXPLqeIVIyO+wVBQsgSMLkFI
RwzZ3ij7RhEsxf9fqYAkjvmOqH4hnUSZhOa+LM6ji+QCDZxgdujOPPvJpBdP+/vV
gTGbbggtjxMtBbqPnWmNCmqIkGcY3OQlF4LjoPrH1mZCkZyoyM/PyrryHrDrFF4Y
KCfDgk0zEWv2I9QGKijtoR+njUPcbety9bkbYU8OcaLQ2WG6uhWJiCAdMc04lfGN
LqfAIBHo8Za3swRZXspMONdKbv7hLhE9EiOUMxlvXJEao49pKLzDh1XKI1Y+kb2f
+mw5H0XXWB1MAK5MwM9IODc24zktkadtXL5EYsPiRSOb63rrvmQNvvJNVk0MeluC
aEALdxo9nSgfWzYMKk1DJgtci3Qw914noDY05B43GMEbXpsi2vB43BgKewEoYGAb
CiVRofi8hhV4FMV4whqWfcEtdMeEIIU5u60mfxmcOaYBauf7Rt2lKdK2yRAaEync
hcBxRw5JPRIIOa+z65fFgroZOTdR++V8DBJpyWuPaX+KcYyBri5txph6Y6lKzkLj
YrW7QKA+4mRvDJmcAJaMKrLEspMGZyPJfaMuBW/NEWXI1KV9iFAzt2f0djlJRZru
vPqqrE2gCjJ22mNA577hYFdCX9S2yHn4uuymQjR0crqlOlk4bDlDTVQubM5Z5cd3
b/sAycUEtFoLvLW+rj94wjc4+mRVmq+BRWf6bAwKYBMxP6XlS9jj0KPC/miuq4eX
uUgqZQyD4D97wHgv+jGZgVkak5gjhRhluGXuW+zDaFWKCvlBnH/6wNb737qTk2oA
RoB4KtwJmOKfaoJAtZ/q9O6N0TX7KJGUXB9osCkmlT2HQ6YXi/QT7ROoTPJdTZ0F
4csg5/aTUqWwXGmUsZ/LJgQ46uBwDvtahmC7jw8cpkyStVq4V/pPJwpNB/mSNAbC
LYUjT1Fku12um3Ux+Q4UdijtAuQ5i7RWmgwiUzOSrmeX4xRfxyLTK7M6EuoQ3bvG
kWu96RyNAH6e35N/BEdOHXboAf4QsIPeXXAXYUyYZovBkcN+hUD1j367Tub2MIsD
IaiP3YwiENS1WrX9otlH5oT5SvNgHMIESRHmaEdFiseUCGVHDV71/rb0F4rRiQAY
BJkb3+5RwOBp9v3vxD2/mnR31CRTVNNXfG7wqvtMz5oRtwxivsmOf0OyltHTwZ1T
q17fWFw0B9ADYAUYtA/X8JRws6EMw0v+zO/O3Yz0IcoMoNx8qKr+eU49A65NJOwj
WpTR3PchorjCD2oNxY5hFnGYroKDA956VdAg60NcEpTsTo2x/GuELFYhbqVSoCTI
yMjiSkMlbrRk4gBTYh2Ou3+RO7Fn3mLvvNORXU2RhRD1pXmRYbM3yklaZGsRrWWr
01Bkujgg3aaFKUXXpOhi9J/85qAwAmMnbntZwdepHDWFRHuT1P5YpSYRLLZlfwdW
BsZsEvprE80TCnFMAyA7jbwlnB/h72WtcX/H21hPKmCTKC71MorJrfjdWeWSzxDq
2mxJ0+PGbc92V6dwVygluOKSPPofk9V+tF24BBAktYZdl6KSqwm2J1uFbda2W/qT
HrGmD/s2IEV8AA1n/VCGwSpAlzSBihYon7kbED2ei5qpZGhmwd3kKxgi2f+x3T+X
HGv4ZX3X4o9hN6jM1ns8aEqH66IeuxbrRZA1C4Prdvxi9ZI40PDwmq3xJ34chol7
7ul82OTSm7bILSLUFbKxwg2tdn5J6YTTap5q8JhcQci4EbGXe6l2wchCvTKIweNI
71WtHnHNTbKGcpgEi8RgJxW0gdwA1aQY7gE10cAnfcYJ1lgL9qDY0JxoDVztIFoi
6jpD44pinU0rwAMy1SfhBT5/iW6OxkioKRSfQeSXuoW3GImqwv0gEXWGNyucPjg7
dkoohV5u7kF/4vI6bnPFg9wfQLp3lpAeA8niV4luEzcFGS6Ean32keEoYydI1/io
L4kbpDx5wSTN+CTFI0jPIW9fkmPCtVLB+P1LsHEfZgoHPqcxSncCtya5/S63ouTI
xVivHcB1gom3sYkMmyRoBLJ1Yxm/rX3JDfTW6d3rbtH/WKzkGU4ew62/27Q2/xEP
yzJUKr9eRzyahyJA5dOEZwnpVLmJIkkIk+1QL66JfX2DQ4xAOWQtYOkCAvrzq6DI
UIYLPHDJXHXMzNy0nwl316zi2pKX99PurxxU5gyqs6xNXtfJWw+QVFn4n5AXo/V/
I6jppUHn9fA3rUE20UPpm/8Ksh8bubrJ3JyC0bUtTDxTi5IJ+FfOG+jQhKbZMAas
K5uVt7JR/gpQSNuk5Lnnxv/y/qjIXTKMwoi9k3QnFBGxTFkyUz+awfVQsWsXw4GA
mniHEa8EZlzGA7zPmLxl8QuFa0ndxV2PmK3QGWRB/hc7q/vy/gja+rA/jc1i+lc8
0qhAySizKnUSqWeujQYB0174oUh1yKYV4GgZ7zHFdv//abgzH2SfDFOWNaHMAb9A
Fnvq0idXaXXqyCpYpICYiW4gAFhqhxIYi8liyJRQXa2VWVr9uHt4eqn4Gdb4Apjv
VWS12Sk30w35rWj+28hlSQivu2OkUYgJkHtY/MeekbroU9229ySf9CF7AmSMbf7L
vOU5boensKUQU8qE6npW76lkKhvEPp0M1PRY7OykBT/6xt9K4eq17JkMFYlfq473
C/ufTh348FgFUyo5GhitERDo1PVn76qniQ6Ku6UpuD1xc39d7Z+szcZycuRm5kK9
5zvHKYj5FCraaBYvp62ZEzx7uaULrv27rYxxMg5iWs6hxv7OUHQedsZNrdCykj9J
y8pgtlyDYYavYUSDa1C2bfoisjtt3Cy8RP+sk2hiEPsW+PsHJnTgGX2Idz0Ogigt
w86JB29S0gCYb3+BMEhVNUpGQf4q2GsnUfhD/tzRiJQktXrSMDr/w0i6nf3jB7OA
nFhq/N3TohcCYkOnx9ZyiLSJ65iRcRvRG8Biy5EYZO4fW6EgmBJ8O2jaOB/rwfA5
EzfiD7dkPdJ8v1+FqOToc7f7DPLIer8WOmqEjMpSLgvbf9q5BuprELKkg3tVm2zS
mBRp4AQ9fJBHRyxQrTazhW+CcWMtSID6EbiTslLxq7JXihFb7yStLz7IET0NMXIt
Ia5ZYzSdbEOnhxXzMjvM+CLTZF6KjjZfKem7x5972k19piv3wU/7wWML1sPz/D0E
JIosQn05E3mkDCVguHE7Ol9B7zo4DyND88ttYySvqhY4NnRXnNUXJwgKu8PXY4cN
wpLNgwoFiI/xDM/agNvXGEKtAG42d4OX+wFdUk/QhTw44Tb/QO4ERPiivu7IN+wo
n7kb8w0FHDIvuHexOCKz4qol2gTCV4iNHOBrbz8z0/e/vdWK1XUmQIu1DhOGUYRR
h6pZqa3bYV+153oG2DtWlqq63nm4U34HZpy+ODiZm/7P7QTVd8kyPJrEEid6Seyx
Hivnl7m5zOap0T3iopZ+Tuvwr1w2sg+Qb69ZK8ns4dg8q/zJunFfPu6JuNDNzuaa
cD3MlBUvmCz1ubcWTxSQRrISqr985bID1docY+BZ1LHYGAPtvqi6z8H4hESH8bbM
EvR9zymlDJPUyVIkACLjbGMThmGcRUwYRALiT6E44pN7WuF7Xbh1l7jnX9D5FwIR
fKaw7q1uH8ZotYrPwqkwF890ITSebii4nkErPOeWyctXPXiAlSjHKFuIN+I6Jgdu
iMXHgU6a9Zxd75ePml0Ifv6QbYvLdon+bXskIqZKNA9RGwW7HYuN/r9paWkxl4p3
YytmFAyV7Xsf6Ikv09Q/Tdm2LzR1zwR51a0h7tGV2WWkWzHPLEGEh51Bh4dsXFZm
FMA72+B/6T8Gdh0TIKnI5eWBzKGzwxdgFrTEu8biNwMuWWOiO1vgpet3fTIG68OL
2Q98thlOCGw99prlQOkVwtfnDkHb9SGRbUNrHvPc9hstk1jN5F/BOXwfZdeGtGI3
1E4pGwlcS9Em9LXXH3qrAkqLEb5XT0zHzOH2hEBKxdlPjRnGnp4iSQeelIovW1iY
h2q5dZIouhYKBiVf4upRZ+WvJde/9GnFnAQUkhU1LxazYcAr4wZIYIdqAZ2Ndimg
yu0fa1R3QfzWInpk19+IazHFDKF5PdCiRUgfj3eW3cnqf7emRoV5tfblQO7SxeA0
A5SDaA/TO3TOU6Q8bZwWWWor8EBCdqKDytg+XJ8bn1pFONvdmYY34uUHiz+ZvNEw
K/XGm1cgJMOWEa8PoQv03BahTwQjVR028OhmrvBo4y/QSlXilxWZk/QV8WoIheSl
nz4HrgxLYoNprWpdIjZuPlx6l4LYPO7BiU+RSLzNGWGA3uNCk6XSWq+e0oK2dIPf
25b9HnLimFSGfBaGIye2XJSR+6o/YxbrlthIKjWINzhcE2z32ziBkBgHV5lxM8OD
YSzeU+toUyqu94aDYHTvGVoSoNRKvsq6UXe+I1vhDskG2RPe25Ji5a7gWmqvhIJX
+3n0VvcL/zS6qHxuLsfAwBKsTmkVPFoh24WCecAPhU+Y3u0uN2//LbqiSgi5u+cz
OOyRAAeMM6s8bwyz7HT5iFVn/a1N4/JKabtJLNi+SHIDtWGuqklKqmGqkjkadbdN
P5offTNWIlNMQjCd9rqZCKwPFCdjXdGBKb/l43ho+5NgpCxRtH6FWRUxw/y/mTX2
zCKi5lVNLxd25jnJ0Bl/ccZpagGv6scavQ65/nW4PCpaLmTpgsZGi7L/yCtCR9jg
Wlrfex2Y1uPl0OWqIUmsk+nRHkDcxLpJ6j/Bk8zBE31OTNrK86F6PrAAKfp1KPWh
DDqlODyjc9AvS86T0EqOQoCqRyQPwpib4WqFzdJO6JG/cxX1q5yV5/vKeBdhVnAA
QZ/2ha7iZF+flWZUCqVf+QC1FS/y3M0Ix4y8vxdUgdK2mELoV0JHWETVlE+5Sn0E
ZLieHzxcv5UUcM3qMyuN8eqv6SS0dKyiyGualSFKi9Z8gOfMM3D/Ubun4RViCKAd
uEBJ3iuRe3X1LbClcu05rFxB4u69o9P7RUVXpKbzGpvETBbIN4zNz954zqJrFB20
hR+80S236oUADGdQMhmVLZ8616b2UNWsGtpOhGduf1ot/VDzd6z7t3J1Qy6oJ+nI
nFL4/Xbmf4PRwY8kKAt7G4HAXBMB15mmVU3clupba9chhPujxNQBpeA1dDyoGEWb
lzXNzts8CQI3I9M1SR2a8vkcJV/9w4DZYCBa9gwQIAGHJifACmZQsPr6d7e5tnSC
jH7QSZ1JDhoA/IfJOPDhn/9TmCsJb0W7qQcgC/dY6FFLfgbtvhbyDo1gFJawBjsR
wB3VR0pttje5lS8/KAGWrHWNwu461fqX0KWL8HGvAm7mQVN93FUwFO62vUqvl/Wv
TaM5ILFNe9Yd/utf/l+5egF6kS48Zta0dcurXa3I2a2Qyhhsa7uprf9e5tFyY/u9
ObvaVG1/ym4jsUKcMGAG+tFU8i9rhuCDYN1HmtNt03vv5Ley2kQsLe1483kvOGyM
T2eRXcCIXl8VNUUNRfAlOtg8Wu5Ag2wPXn89801HGBEy5ffj1bA3Q14XuqPUHwvP
iV49z3n5d7vdhTUsXYp+aj5FekxIkb2FC0P9xmWmGwkiQHzGNsGesEAU3TX1hQTg
3hgpyCcRuriE4jT6JKTDfOTQn3L3BPwZvbZ1T6vmOknxWSz4UY75CnytZwZMAREu
UTSZJPUsd+5oyqyFzbeyeIZg0r1hdA6LKM3HiXy0cpBCBbz9dGpgUg55Pe/fyBgW
c4nE9cCgMaFZdk1tIyvstkaPlDjbs5ishBuJQ6Xb1NsyPYix615Wlh82zICCtAXG
3o1Tp7c32Nlzdl6lCUco/jIPBb9zEnJGyh3j9N8/udCC90cCux2tU3K8xemymBWi
Qe/ytjhBO624K5efh8aVttTjphSPNEbCU4uTHrFORRdw4dtDE6MYMJ23/HYlGp+O
ajsJpkkbHMP5QTl+1vjtm3g3USVuL1yRA0dplrh8oU7AtHe/SQl17C+PNWxHMRMi
h69AHcUt2GJMTAixZVY+3vUYzVDU/oLyMVC5WW0H0zOm/osWXAOEhjiafTFxLbC/
B78uIdUoSCa0B5ryB8pVRYItLn9XLapkpE/ybGmPgjsHSTR8vtJT/3Ev9vnNeviW
IunxY4+wN9lDWA8MVIxEi8U0khydhw0PSnCBGD4mWKbq8xrEJ01F0TknmHwrAOti
GDbGqbf2K4VIarMQS45VqG4GTnWUk1j80QB0ndgvf1OXKId6/KSkb1WbtLCnVPz0
jYDcwtt9DHzXk8Waxqk+oFP+HtAQvYHcVBbMJsEj0aj9Ykap1wo2bI7OV6EEOlVd
UFvZpvqCuuGIFvWokXVZkFP2ZjKF5DAAWkuhlpIQeuNjQ2Um0UVkSS7xq02nRzJT
jBTJaVLH/XFCpWrMXWju6HAlKETE76tbUVodIEYKkN81NEHMJz+AnCDi0YoYcKN3
W6NBLDp4h5FB5tM2G850z6x09CCqXIbKSzSCjcAIhwFx3BtoTpEiPvJYuHILw3GE
kFb+TKgl5r9nWmbMYx8+kz4afIIkBavYWgOnw5ZOYwQychsTYeNp0yspRuml29IZ
xJkunGqzGyvQX+B8n6dXtll+mE01SJDckSmFUiHA80rKnhKiEmydUZk3u13wndQH
KOyoWtexAZJNYyfbQ4ZPXOT5W/B7LhHENwEISYi0ojWuiMmreivtV3QbV+alof6J
pC66NR6m9cUzQpZc54FIxy5nBcv3ta5drxHN3KFI4sQaUHRK6MLSEbH+mhdl3TvO
fLHEXVS2Vjc84ddRo2p4F1PS/r9LFHABNjn6uTRV74/uDU2SjU0ngvXIigSzitU2
ohjXOeN31j2889WGdccRQFZv7tt7uFezbEO6wXNFdUEGFpJ16VLYVVi+QH7EM24L
AOdjmgs/rtkxe3AAaei//YJ+rqp0wicbuflQzSXECfI9O6Z1gNYENSmha0CXWNgx
dZdcK2F7C7AuZ4WdqBG65jjEsjJUe7ZLAY12YoBjxuM9M9KhpbLkDGDZFs1KpWe3
vanIgPjHTdtcyN/bRJ2B7Ss7nT6XnW52V7ZyVUrpUA94T7ispE1+avp6qeH9qrzX
UC2UqK4287IlZ6IUtx3ojmfjINc2h0n6xvGqJ/qHxjW3s6JBxY+v3US16OVPeVYa
jkp+o3xO0uQXMXEW3FzaFJC5RDB8i9HtMvPoym/Fxgt5/P80ggc3AzKA2MGUURYP
MfPgCFx2LZ814j8xBCjjIgYUHZ/A6GHQWwctflRTA39eDrUsm1Gup0y2No9U0hIf
8rkPsBK3SW/IC7I1A95FfmG0jYI2gfmaRS52uT84h8BKsShLxbjPluZ+Vtjr1F9e
WnRa8sjT4C8ZSQdDJklJE5zHVRxXDKMGzZkgIufXUCc4R0qwJQyMyN3d+H6m46DD
`pragma protect end_protected
