// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:52 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
IUWMi+48xMJgVvJem8Shg1kvIf5NenzfbNPfAqLDI7sw74Afsds1k+57yupl5ITT
eFpU0ns0xq9hK6XoizbpgteVEOo8S4ZBhu7pzxT3x1vRrzCkWb1dIs7qzrmFgzsx
CozDBz6mf8fI+35IuqzSgOEFCcb1JqQvBjcD4GtzeeU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2496)
AOtz6SZAAkHSb6rPliTKv1CR7vfkPe4ht7HwauhUl87TY6Tnl6VF16S0fiQ1nmhJ
dbW2zKjEvXV9gJHMufd9qtuhltqgIBA5yxprrTuak1q0mVxo9qutkDumW3L1sSc5
Mh4cjiI826xBG8no78V2iWXpwoJsFibCqRUVh561wN9fjZJnaCHdYEP/0V3Kxnj7
eVb03/fNigCDoeurnul4kkVZEa6wxUyhuu8K0Zd7Dhfrl40AUna7XmmvY2vAaKtY
6K+oLg5EoFVHxU/KPPWEBVd+iy1g5gc41KbAWkc4mGc6ceYqljVKBcuQ4oO8ECIh
VU+l5RbZUdJwk+HjAZtDqIiXG00ynU/n6JgwsUz2KwdAOa61LY/BF2cmiHpsATPA
hZSlYk6eTMyv8vOxLolNVDhkeQgVSIfgV+fgeJmJUh/gNNeMzDDgMPDr9lnsl1c8
7/ydHabRFUYwqXmSjaaNJ50R/3LNVqIlB/hmiNJVgL1A6nSD++zpLkSiKk4Wn+NJ
zYlOZDjfVW9pbkL5CqLnab+j041GdbwUyF5OOLW5djvKMD28WpbLz/1MXVV+EMYV
ZZiWYJq5WS+tYlpXI33SOzRCROtlMtp96dIaaGVg98tGRU1Aa1MRBCI+eYuEHv1+
qDMWUtliFaxHGrVX+ZZjIaepxTZhCQXAXFKRdI5ruuAIe4ohZBv5jygSJBI/jdpO
nKbLxnrQTS+RFz8Jqm7pwMgdRj21HUUlCYP64Dhj6EEU8Z0ipZbgKKYAdSc01oMl
3NB2jq/5Zg5FUgwq3XzEKxPURxDOMME9JxE9Vauc+X/zPQK2m9ETtjs0M9A/t9q8
AKGP5vatAQKRaN6nBUiUd/PrFOxq2HFb3U3mKFYjf33+516qSP3qLrG3NnVPsOlM
YrQLD9aRLPjdISnrNKQy1Nf8+ZTLDhw3NlNigTSKRs3Ez7JTdAJ62QAU1jPEto20
Ceg5678eLBciXlIS/VjVp8yxLnK5T0xC9qurWTaFh/6xWwiQLciEED1WJS8eGaZs
TKW9SE7PWkL73T+Qnwc4UJ+4HhoKiatJ9EfXpTe/2x8pe/7osd4AhErh8va3CeHr
wHFyOl5u7K0DHA5MQg5Azv9q7maA7gCRWNaIfN9IQMkjXu5M0OBPTJWJPjZgP8KU
paHJIktjv+1DEPnc9LDU7Dx0kWSfXO9J1R7he/s0JaNESgVA26Qu/4uKgb690dpk
YFN9+ur1eATMl201QICZ8gEjIwYmyk4Frm1Q5eZ8tECU/Ppl6sAh/etmQo2Z+rAr
garA0rzymKnX0sRSJ8XQi3JHncAEcy5iC0Am1J+Sfs67k6aOvseOxp6AXcuwm9F0
qy7/icMv73+39/UTe0q06C2SyQJwXxCvRp6y+7+cS4l7bECyLqk6hW3PNu3D7asB
ILHB5b44PRPk8QJKmNzmgFjBIpiAvxswbSVeBjiukpc2pGwYklW3MbOdMrw0oSKM
EHsiMwegro5EohUm88Wz7a/tGD7X+hNxY7OXHSjz5ryWigdJ0ytUGX0vvmbXU2ar
BRCT18szNelYXtpIFkD6EMdhcZHeF7hsqVu0hfd2rl2Je1yqaQ4ShbxbYjPuQbiG
efgrX2UlqaUren+eLvBuZZNb2HuBcSsJvdpf3eyNd9dqiAkyxdeiHlWJOkydcUmn
l4B9pv3whg8Z3IC72OZhodnyHXA9qKi0lU7soLKHRmF8/fFI0RgPwTLF3poKzT2w
F/eJgUNR8l3bPSNmvavm3boH29VU2elPZaakSUJs05zxYflAKGEDliC82Va0os1+
OnihhYh024yO3vtckI7uKyvUGPbgxOzAITKb0Ftp9B2JxigwoxLTu2AWoLjySdlJ
KqDtQShjEvmdK5ICl2W9i/YKmd1OT/hALZVJdgFRBErc9+jznz8lhiIaDWT74PJa
k1TXzc75cfmSU0WdF7z+r90FWNXgj/tqad+Xx+Ay7wZIzi3uEBI3Cs62LRc/oUFk
cqMiehgr5hduGZXOWA8HNgjdBC3uEgNZf4H5XPP3kzyvEbsN9lPn0pvnfA3id0pE
wwsKzb0Os4/Y0D0imPKXZpAkFO0Y8bajgc1XMGf61EeAibG7R7TXinkM1x7npQPD
N/16eW46hcGAqaU8D67PI9dmE2oaOTvhaz7wG7YraUTORsHeVP908iouyJJaMFon
j5NWU2ypu1ejmf+EDnuPzI4/RIfK32EE8s18SdTpV9Rf+gJ3r23P0dXfC0Pd/4eN
tAGbEPDY2EwsHVxH1XocOwDWDVPoz7jDkJ+9WkP8HZr7QbsnoxqcKjQd2z9IDo+c
jziFa7zdzxnYHrDigj6geHHb28HGG+awd94C18cRbH23hUOMQUge74QryJo5U7Jv
r6saA8KoCohJLsVOrj2MLcQmpJmUuVlj6JlN3zsD8Ywj6ESZWV3WtJXGT8ZgM/iF
mDdkfZjc3bP7ho38WuqZfOt9s/bj4RES2HXuhmOHH6ThJyLDNFxllLUn8si+ZRqD
NGmu2TtcnAjhlJfeeF5v+N3psnJuPaLGr4yr2cs+S+RwuRRq3nsy8QELuCsZc64S
ALUMCQCZ6UpBTLXmF0dnj2oGtoEaOOx+6/E8PHmGfCq4uHS1N/zwPCgt0/z2ZoeI
NDuTn+8yUCd+/NF3h7FtoWRfvK7mwYNF9otrACV4zQbQC4b+aJf6PrYYlJDvEk3w
HAm3C8KD+v3oe+oOK79QoGQrrMH2LgSI6eperArLLgkKr+n+z4S+17F0yRHiTmvq
JQQbnD6dm/rk/vNtmfoXcMArKYdOa1PTKsf4gEtngJsGd+feZMv1d/HNBulnx4E8
f6oBKJ93aqLzfZIXIVxnXj3RsHhqhwnEzkyBNr1VVjYUsgylgKFn2WpBJIrfNL6s
/dmyyXQSeMCdzRV3GUXVBB15TvBkpEvAU34TVlpRe1JB9LN9T+lrglBfDILAlL+V
iv7asA9C/PuD2o5Iig35RQCdzLRIIfJGVWMaqH22nXX3T6g+9XKNsInSnhh1oL0s
8dpJmo40HLpgA7goZJ5qOWX5Px6bMIiGCIQrbBstStgt8DJO2J7aLeUtgR8cmj1+
Dm4uxcAv2V34VtX+rsBApIPdstSSX9DXv29qCAIKvuhBMmJQRu8bNffAGl5n0n9i
wqogxHs1KbXHr2bNJMOl97YRLdR82/ZkI5TQ/7eZtq2yKd3QgdgPSlXU+BTIGqny
xkCHJ4H6r951CKNOecoeBnlN+zbwzytNyE7cJoq9mGFWTBW95RDJSHaDdI0hbq+m
+CodZsl+1+v1SqyJ2+MLRxEcXQdenMggsZ4Qm+ECQammJjSCwtg3j6Fb9zVf+ASy
`pragma protect end_protected
