// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
`pragma protect begin_protected
`pragma protect author="Altera"
`pragma protect key_keyowner="VCS"
`pragma protect key_keyname="VCS001"
`pragma protect key_method="VCS003"
`pragma protect encoding=(enctype="uuencode",bytes=200         )
`pragma protect key_block
H_0,Q"!C,; 4,DP4CKSQH \4:</92';<(+I6?LP/M8M,$CC)"VQ7Y$0  
HD4U-QP6U]TGM^^6N3DNU!LHM!7(W=3[)?"><VC/HD^[E%PXK?N? 4   
H<Z&V\3+A)47R<V)M7.,<$F?/L:*0::G\; &#G$UR9(("R#LYVB,C30  
H[S/7YRA&S$G@>4ABH#+H/ &M5"F2E_X8GPZ'1$D99^-:Q:(&1:\*/P  
H!Y[+U91.Z)HZ7CM\7:[37]H<1EOD>O_@'=?X5]X6*1?6W7.<=_0OL   
`pragma protect encoding=(enctype="uuencode",bytes=18800       )
`pragma protect data_method="aes128-cbc"
`pragma protect data_block
@S?)E=S-HHV#AI]"<\_D*>*SESKGTP$R2J)N>-Q_)+KL 
@#^XF!D%*):IQA9%OXY).< UF=UEOM!T<)N^R>4)G=\P 
@RN2&1)EX5+M)_$6P)+[)!9N NLS;?P4T-7WH_IJ+988 
@EO&(7PLW]FZVZJ8Z+W>8.:Q@X=D,UP0.YN7V%?_1*ED 
@1:FC@\A!D;>#)$V+K D;\LH\GFT^^KOGLOX[M*-=N<8 
@OLC)<Z 0PP5MLKW(?(E!Y%9BK@U8;W>.(2G7LM5S^), 
@@4W/X C-3]*6GJ[]V/JU)57J7H*I2M!B\TY.%401\6< 
@P8F ZN$+G,T$.FH/^"KK,\[8_X#=,"OOH".$5_N8?=D 
@LLA9S1N8LQ?"L#-1.^Y5M)8]MWM#/ZX6WHF3SMI".Z@ 
@ RY!SMXY%!^Y79)1#@1:,)%%0%]+ !##AQF^WY,L76, 
@BE!*LX+S-_PFS\$FIN:+\XYR<&CC-&$)%:S"7PWK20D 
@2S\\P;VV0349Y6XEDG::>Q$X- 17FT<S.*I/ N!?:?0 
@(YOJR4 506+@(\'XC<38&CAC/@P<#M_?YYG1V *"!W@ 
@\$B9WW^L,%C/\KK"-N_8%757U6P5'BQG8(G0JE0Z"BP 
@LR1*D?<">_4_T!(L^Q$=<37"&I]ST)&\<AO1+<A1>F< 
@QO5Q-?VV6Y[;W4\X:-C@[-(U+J.I\!/:E3]Q$$:[KYD 
@]#J&ANL-ON*-N/O'\V+TQH-9'6G2+(D9V%(7,IQP'], 
@MSEMVGXOT;G-(='SBK8=Z/AW0JSS0EW&;T]B@O FE$H 
@?.M/Z_0G=AO"@U,W#&4(-A52S2\(C9$7^I [^51')'  
@MZP5/ AWVYOK%[&C32UL\R5!(J<WA'Q13PYTP$Y>M=L 
@5)P+SD[I @L&B+M\ O;M*7D4(S4XHE\5 ?*GIR&E)-$ 
@&)(X+%@Q4<O-K\F\&,8"4"YDW!3>XR7OV1M%8U_HCGP 
@#TAM<RRTJTN=U]4IZG WG=3P2\-^0Z_U& D %KL?EB$ 
@5G>=$OW7@W[&8O1HQO0PG?_4PK??2<%$.*'1#P_RUS  
@A(AY*KW*\RR93@0&+=0@S!II*^TF07%H5\?A/?QH090 
@_N;-V!5V?+8K!X<S<99]B(ML:EJNBI:(8:=N4ZZ3]-@ 
@"WS;DV9-WWS>X6BC/ ")?&:^P^L8D/AY0LAH "D&7BL 
@DV9\_ ^ "G&9.ZUY&*G"2?0S%R20KDZJ07:0GWJB;.0 
@K80ZJB'UA:%EW<<#A.H3;)XR<SD9H (:=PT9YB8P.AL 
@-N>( ?1#\!-$:5)SRGCZ70:QLS,X_),%-1-0$PX\,P8 
@S=O9LT*%^<FE$6N&2Y.906J3G=[4C^@>P%1(@]8^$KL 
@44M4)N#F3C%SN(5*Y-Z%U*-+IE5,Q!D@F"2E4#STJC< 
@8A%LKWB1'@BD.#LIH"\ZA/=.=5MU;WI!(-38/$3\A>D 
@JD1G6+8NI?!K _LX9K$>&KC 8[&&']YIW'AN.])K&V, 
@H-VO<A=G[:+Z6/68:B .SGM*7S5<B6?P$C(-=DNV+7$ 
@C7EBYF'J77:X;L@[1/00FA/U'C2O<5,!]]:_(ECYKG@ 
@5< "H]6AU [+ VD&)9<\1VM!OT(% '3#0?XI>H3ZQJ$ 
@3L[<BX4EF_YUXGPQ/V7,6/PT![R>4&(8@CVD'&3W#T( 
@7R"&!_JYF'BZ[22"K\=C;B\'Y'8J"1@MS8\-[+!=0U4 
@^F+)/ /6K8%:D(L'5>*!:HI<:QGNF)!V2R!J%H*)ZF( 
@<27(4]]PBI%_'$9Y9!.4.Y"/0C_ QLD9:1KYTDEA@C( 
@A6<IA8*.62U4:#]\N>Z6AP>$\EXVADP,J:CQS%)PHNH 
@YA@;<XV7@Q>J':<@2ZGZIU3@P0B"Q&\-M)$9@WVZMDX 
@@COI-7G'EJU*Z"N^<$[M6,/M8P.^,%NC MBS%#._S-( 
@G#<WNI&^G&NM7QI+(W4:+C_;$G44WK7W_0'U<#8R!UH 
@N?F@6?PEES.KTXQ"S8_7F[*PS#K"IG;TC SX6N><ZOL 
@18<WD[D*")!8?WMFQ^?$ E*Y!H6#6**/#*+]VP!DG;, 
@0=0#9CTM$?1MX][DF48? RCE04WI4OD5HOUXFT+G]=4 
@N%/%"*D VB7U/(E1HB:4,"HC4:E[ELX<:^*O94#WE 8 
@2=X%<UG<>'K><V-*7Q/93BW#2&MXI!-^C(J*C\+0"SX 
@'IG'WD[=A'I_\'D#7%70ZVH&(+\=CDU6R7V  1#,=(  
@7\Y@9?T_R3PF1<B46VX/_ORSGL1"9;OS*7-<N/E($ 0 
@VIUVU$ZQ>54EK>V1]SK83]B@?)Q:8NIV?E'A>,LQ6)P 
@S^,FQ4,D9]UP<6L;P%) AX!]V[B8CU.;K!9OCX@SOI( 
@630^,IXW0.7& T2CR,7@UZ /Q&V@T0_6W)GQ%F& KH< 
@-*S@0',?_C;;U2ME1:)GA@)KJ;Z?G:+-1KJBQOQM<QH 
@/41OYK#R?9%=;VRDTB]N232"9Z8\Y()BZG#3G:]P]<L 
@474OEP4YY6:T="GO9 KT(LWS"5I%=B)9,$(D\MAI*1\ 
@2:(9I/2Q[K[%>M?=5*A. 8*Z5,;84T\52(PZOG&+;Z\ 
@E5[4[<M@Y\M\!$G!DU9Y]Q#L_!<J<T79GM(2RAV))$T 
@-UE8&V,/;C"QE89T':KO'&8W0M 6IMD PCX:HTWA-(X 
@[CIE*ZU$"EY_@:=A[HJX"^T@ZF>]?;ML*;>,0K_W.+8 
@&XO4ET9Z?.L]+,B9!Q@_X8$Z/1IB/\AR3]AIQJQ @48 
@G4L5"G3-G9YH&DWV[PMUM,1;RP'PE*T#-PY[BS6<1)L 
@.>,JH-D:.9Z&?':@5\$@#]"@ *Q-K@<GJ ?YNJH#V8L 
@,9WJEW(L=1)J+^LF2_\&?24QX:,W]2MLZ>" 0!O70.T 
@L[,&?ZQ]GB-2'P<3*&[J C>)CY>DYJ:SFI4+N;R%,9< 
@%CC&A%/V+UQ9[^FU4RZ[K2#RZH2O7&CL-^1\*U362B< 
@9\I]XZW8N?,.MI?<$SIPMO9@@"$BR3%!94Y ! ,]67@ 
@^C;#KA>@GI'6_P]E=JXY?-VD($#!;_3"M'?<$"(21$L 
@V)OK%J>2OI%S\^4;)0UAEZVQ])!Z8 N*<]/M>J?C^@0 
@3E^RPKL+KVKPBQ]-[D-1 J(+O7GJ5:(4=:Z3VW5]8B4 
@K5!H#>8B7-_SQS95QQ%E'GI-!.1^+V S2&.E5N'AWSP 
@-4I$*2V\VQJ>'C5RPU47&!G)K(3(3M>G'M:OA,"=(\\ 
@_MS$CXTQVC^OPTYB$V5$=8@I$$Z)F("*^\I@@6:][Y@ 
@%:-N&M]=%D*_X%G:NZV#IC8_H(GRCG@+5\0P^"U^6G0 
@6^_T;V\BH)D(CJV$P3O5R1_XI'6S2#H !CV_O%O,F,8 
@QM T .?%6MYFG?V. O.T+O-14HX&9]K,Z>CE!+1F?UT 
@2EV0NXKG/!#W:^&/ZV42'O? 0CE>V_(9QMYFB/]-KZ@ 
@](.S8U>RZ'*@#<GMT&*'?!X'32P1!FWXZ/1;.3J4"%@ 
@&'3%2F,H.]'+)4<^2HQ ^.W:I(=]$Y(Z\ACED9^='9, 
@G\8T#!)ZL(G&M.>>.8:_S;CO/H_GA9++E&T[&.?=CP4 
@XF)?]/P&O")YGE##<Z6#?5AX?8_)C-X0UX>P2'&HDKP 
@WQ63)SS,74S;!]HK$>MK4Z"-&(%I&QXY^L >-*U%PP$ 
@AV:W,MSJGE3SQN0KQWRSL UC@,^D;81+9X1GGJAWZ4@ 
@0"B[ETI@&CR1C3ZCM]*0NF/DXHZ]M,1>@'S!'CU3U94 
@2R)00>!%@8PYN$$O:TI8C)*01#+E&0(XN#R-(./N!3P 
@#6RX@Q05IA"\GC>U0Q)Z72$U:^ := IP".U)@C HPX0 
@,_=)%Z)[VXA\"#CR6=[YM<DCE>0Y2RJ$11XM1"&((<( 
@X./IB4#UW)NW?Z?VR<I-;. #.;"N6@,0-5C4R,;2(SP 
@@6D5#](N!#RU (_LQGCZ(D 0X)0ZHWXPDXA[L?!!1C4 
@Q !AGL&5J]>#YUQ/]4\OU5O%B^V& ;%L'[RJ"U/<]E, 
@$IX@J1^R\4,&_]"(9ZUX' G^W56I<EE8?%J\#\ODS%0 
@@EGV=X&1:&Q-9<G7#Y+3-B-.:K)\_"F*$XK/GVJ8)/8 
@(GY3FF%EWH\K*4VEKED#(:,6])).K:T\:)Y4<B^298L 
@9Y>64&:SB:9\4%$#;:UA@>*!;PIM$T%I'#3U_>Z\;&X 
@+;+P*GIMZPQ<.XF:EA_OQ]9"+IE.">I2X)JJ J*C.9, 
@&S5VW7\$1'LA4[0W]+&TS=Y;!L*SD%S1:Q-MP&)6KZ0 
@J3TN[&+$Y8.G!I9O1HZI@K+-/"8_K"B0-AHT16$Z[X8 
@L5@9=E/F#=M'T+1I=DV@ ZV[ ,0J=8 8XV\ACV""($T 
@_T/:36MQRM06"F>D$LT1768?@RHOJ\\]>P)B+X(=[S8 
@S1+"3T DZ'GHR*I6*(#8O9G\P*X8?SXOICA,QG/__C$ 
@,;%]'64=Z:'_GG3:\)(0RLQH3I"*-PL:7I 2]3[I0.8 
@A&((4D6D#L)F:( <COY@HN4ZSV:3)?TZCP@MLN;RV/0 
@IMRS)8+SG8DX";DZ1I$H>KH4R?'1L.2.?0<N%TM0?QH 
@'T6;C'G%"%U"1\C3=4J3Y%/_%_#E<W9!0(<7)P@]IL4 
@IMQ,@J;#:,^^Y1W"P[+)H^S^1*@172F;NW&:#U$GWOT 
@%$D6VI>W!9SER #0#,D>8<4=-SG//F8N@OGJWS@BGFP 
@*6<XVK<T4V8[?03^Y@FVK=N0D<UI<=:+U$G?-FPP[=8 
@?Q>-+V11[ZKFB13H^T> -WF4XO$7YO1*]NS2HV/(5\4 
@D)M8&+70R]##3E"8LU!$:$;09^GWD($=W6FI%V7EC"X 
@QWF(L&SM9%FG@@JUBUB@*6%RYB/YV9$00#R209<$P(8 
@-&L$"C[5]%\C3<RS9!SR^T/UDC8E\M@XBF3'I!8G1LP 
@6CR!@_'>GW]K,<?+V"MHQ-+,K#D-UD8$4/G@YPTVFU4 
@OD&DGJ.//[ER"V["]37?LH83IE:?+4TFW'K_D,6C<P$ 
@U /QMCU/M!9L-[,,9LG,'W ;AA2')2[V*BX4<C)GS], 
@:K;A8@/+Y?(BP*R,W ?^FTPZ=!47!"E1Z4,-3U_J!2\ 
@;>U=/ .P]!^=-5Z&?,<9(7"DV)(]\,UYK2*,!9OV"UT 
@Z2/#-Y!.QC? 1 P--"N-Z,AYS?\R1'[!P/V0IZ+]G&, 
@FS+2GM'T?O#,&+!(.BQGH6X9 6QV4W<GAN;J1"&VF&( 
@=44W)KD/$0&OOB2S_2J<ER;M$:6&>Z6#O/YF6J1"_0P 
@_Q-6ZMD8 1OI22Z=4"-&Z[+0@*(MSD#*P 5#.)-5WYP 
@6>!#?*LK6$HN\IME#2GL2!$0A]V/?NA:7V\M++N5 :D 
@XGZJSJ"Z-S Y$G1XXVV,XKO?K!;^[&++"4/5R#0S'8X 
@X7H'%+FV?M$=DMLTL(E*[.U1QX&F_YW8-9T;Y>?=^G, 
@.??^-S^LTC@[Z/[)S,*D4$O^$8VZXH6#L.;7[ELABCP 
@B\M]VVZ-*MC-<=#]XPO/]&$'!WSV""<]]H+W%[;U^T@ 
@.[&20BVJDLYWMR, ;:41K$VAG/-U]9,]'R<*8 8,%"< 
@Q3)[!&A*O#V[O3#9+>8AA Y1UT(HXWZLSN6\,P;FC&T 
@\Z:-EY]EKG1U-D8N(U0)^Z(AAC<5U*[*1(7->".C%^< 
@FM>(V.MQ%"/=.VG(?/_KH;D8I]>U:7W>5U&6=1B!4]@ 
@?"&;=$<9OZH4'H?V_WM,_8L_I']?J0D##S0L=S7_I&< 
@]$FMHJT>Y132/S#B;C OT:EY[2CNIM@>F;#Q)8J&G$T 
@/%E@H27+Q>!M+H@>(,D;BF8^V>%4;C=]_:36;-V4H1, 
@0XLSR88O8H&*:/%,ZXAH+=*%(7\:.ENXT[B!^2CPHL  
@AS5QOPJX/3#.&N;NXA70Y&2X)_+A(' -WMC2<IN6#,P 
@^GY8/PXR9_I,8.&FVO9/3U *,1/>FQ!25T-[]BTFVS< 
@#HWD[0:#J<B>:3X127AS)UOPV*N<V+S=.%JQB[)U:N\ 
@^\/??83N>N8]B,]F@3Y/F %]L^.[:T[(1MM."?2+K%P 
@_/$L/J!**")@-K$YR]\+4^'M,*LHE3,HYY:U7]JD5Z, 
@W8UGY02G!?Q.3$J9,;.>2\M(RZ6,;5U#@VL&YKB1>*4 
@[JC'3V^.D7U"I]A.R %IE=Y11SR$LK&E29%G&/OP-/\ 
@ I8]+>]L^1>^:<,.N*BFR>JJ%X[YG2I90%8V12;=J2\ 
@M<%WC'+W[ -KH WG^-[;YM+41$3!FD/CYQ&X\EW>70L 
@MX 57K0)(09SMGOF;FN5_R*9A0OT67KOY%U<Y$GSY7D 
@5EGV2\.3\+:6Z7&0,Z[=@*J#R6RPBY3J4YU86+YX#PT 
@F* 9]2-T:$=;LG!F$3!  O2&FH8BY%H7>SLMTBA&\)D 
@Y:/%!VI'$0[F4@?%@(TN)5/S-,>\N%!:^,=F;F4\G/H 
@R<00G!$VJ$C;J;C+FJV7MI'KZ8PBK5\M2,R^FT^O02P 
@BW)DE>@[_L[W$;AA8 =$SD16HF]FNFE%7WD/?_"?  8 
@I!3M-2Y8?[Y@Y4?K=1'\I*A6=F.\I/9V\39K=)?HL:0 
@K1E&M,O 9^8"/-F7IH41.I3@N2"0[Y T8@(^,7;G/+$ 
@M%:\LHTQ7+=\.F+X6/V 5J,;#530!$JML&[V%/3?AD$ 
@,%6WGQRQ_,[."%$I",E[>\8ZU&31EKQ&$M[%4S]?] L 
@?H)L2V1K""*Q2.=!N-C#^H\+ZZ:5+LWO7QVY0DT<):$ 
@#-,:145CR_.D+@_<?HG?UDX8^;/ #A^W7/<?SCE 5:4 
@E(H?;T.=^/7S6P<N0XTV0 QZ@#JD<$>IB%?<6Q(AD14 
@4WU%YP7,-IED_/1XU"<8DCQ%/;'9NTXL+IDCW?$P^@$ 
@D0_"\'H"SR>>/H*<6H,+I<"D 1OSCB&<H6.>,.U\%HX 
@14+49C<[7Y3Z;5WBTK?< ] !*G7S2<!4_UX_3"[,VF@ 
@?JIE8H< @: ^/]UOB@,\<S7A"OJXWE*K2EI:.90Q,C0 
@+VH+C/,<_^I+1S$%B%XYL$*P/2N\:_^=R')+VZZA4N4 
@78\PXH\0.XRO*1_^1A:7L\6@0O1',W#P^EQ![;W?F!( 
@)3^5 1R[H;HWIG[IEY775(B,CC1V5!VUU)DX\X#YU+\ 
@%K%Q=:]B31X]&;(T!7N<R7D("%>PG>'K\GSG4&Y%W,D 
@$)VO!]YI08$@,-=F9E;5V0S_BN(&M+(A<MX46FV?P[P 
@Y088CH<(^YGCQ(ZDCKB;W3$04:QNP1 BX@N,B5Q.+AD 
@&] U*79Q$(?\+C!;ZJ89YO-:$EN(EU_%E3[XTPR/[,, 
@/%VD&<E/A[Q,?P^AB"OM(UJV24Q@ +K0(&W*2PJ_8%\ 
@XH9T$E<J672210#DGD%_ P6Q)OU"@3W7@YE5<6&"[^@ 
@2O=U0*<! .HX_I3V8XI:!ZD><Y<YV<?BC,T2HGF%E0\ 
@0EEIZ(OWGR \.U6#9)PX7^.X*<>5-LJY.D>T03\.UZ8 
@O:WY6Q4B3]@2E%4Z&NI*Q8I ]H98[HZ-7]_QB'MUOIP 
@X_:7>G/RFL:4I\Q2'$2DM0G&AC?P.(X%%+<E0BGW(), 
@\"VSBAB9."T'@D6#:J5_.MKN!F> ]%JL(-Q_MP^*Y04 
@%BU]27\D  1J4S&]GDER!:X_-4%Z<%O*:,3,1[J0XEP 
@1NG6 __>]_0\5-+O@L(*X*1KUHB#.'V S3]:'JZI)RX 
@08?B0[Q/GQE#R9'RHWI?=ACR)]\S/K!ARAI0OA24XT$ 
@(6;&AQ7KA_@P-_I<:=X^0&_O$.?SLV8I^KQ<'M2;]98 
@2Z_O^C*%_L6_7E8KYJ1EKL'% S)'$LK#FWGLCE)!1JT 
@]25Q9V#*"<Z\:?NU#+ORI2;7.;AO=7'/2[#"@)AP5[0 
@=VIRGI.8.B#]-BHW42M-BI6$VU^0"@*8"'H[J!,LF.L 
@I*Y/?@[=K*1;0E*$+I9X5L 3P8XT]X/C,)[@;PN-<"$ 
@^=2C%6]Z&R,Y"-O9A0*"5VXZJ"KH2NDFXHVTZPMF U  
@G<I13<Y3OF>FBNTY)\8@"DKM"I"T+-I;\\*-OFT]6PL 
@I#^=Y_7+H89YWH'A=V3W*)&P=6)FA>>YJX=HJZUI)%L 
@OWPD11Z??"7VA<G&.5<O/V^.5X7E+N.VA=F*LQ)RC!\ 
@=]]6=L,&CB=273I\KP^/O63<+R-/_(IHRR(Q2#WQ)?P 
@8;1F\59"/B=:K41/^VGF=!/9LA.O2K#2*4E-D'C["80 
@';IY + ";K;(ZF;TS?W$!S]$&?H<%[79X(4>%-_DU?T 
@29@,JI2H6+-\0&<&#'ZO-;JW_RIF:3SOS?P]W)$5)*8 
@U\9)NNP>$0TTSG6?T'Z%+4O7_;+G$8\,9;;EGT7J5)@ 
@(_+W?X*L^.("0"^>HG>!;4@W0K&SJJ3E-@=\FH5JC2P 
@J]N7:""2(*] 3,'S3\=^*%FF_J"M\=W^YSR&-["LR2@ 
@9M;AIVE*TB2)?O4?6(35P&ZO,)PZ:5I>SL,Z,^W7!PD 
@.NS$)KS*/@X-4G4Z):JS 10J1LY#<:=]1#Q,LIP4CR\ 
@O2#?+8P PL <=C:Z6P!<6SL4/] !V"/%L!,/%4WO_6@ 
@!EO=.P)CW9W/G%9"#;^^\7CN?Z%N/G.V4SCB&351'F8 
@G32'+&;EN\XX90AR0--(>Q-=B%%/J1/.=-]J[.%GE@D 
@):/Z+_IB<B/N?2-!I;Q3ULNCNW")C(C%UH1C1\?P53T 
@D4B$#S:=,5?T"8E9[(ODZ(D?AZ#TT1H[XZKZX8QWCMT 
@VT=-W#V#.X&RZK!9,-A"81K^>>.4&M#N=( 9V@3-Y$@ 
@/D:#D2(K\T\GS'W9):0TN8=O"G]S1>6AWK3]:'%OQO8 
@[G@Z[2I[Q,*^$UD%/^(4Y!()25?4MH\57QL(,K!OH[8 
@K[UW.*H^(/6C:"'"=/A$>AU[,X1J C^V/Z&.7ITS:BX 
@?#!A'C1*GS:2VID0\@G3I)[+^-7,S"QU1\:IQ&K*[H$ 
@H>7?;Y*8KW%GV97B1_KE8EL,M J(O";'?/VIYG_L,4( 
@?YILV"$$E[;R'K!'J3:J%-4X=9.WEP(A]U2L+:F<7^0 
@)"TZR8G%<VVI#+/29X&(^:(Q1;H$Q!L&.G%]E[4VZ[< 
@W0X%"KOWB \^L;C;,2]K"5C<%86SUDTX OT/W_4!\[4 
@Q: -3,)[.5MD5RRF2W</4#T=:ZOT X4N&BZ9@'64!0@ 
@]SR3@DNY0T2E2M2+K]D5+MMIB@$$&>,M(>LK96M,N0\ 
@!%1_#*U+-[6R>J&EA[MDKK6Z<+HM%X-H^4:;<^N@>34 
@7MKMW$4 2?-]$&!SV7F$Q0,W4;EP@,[/' ] L7(,<7\ 
@EFJCL!^L#5EJ>HO_2#XZ^;1G?$66W]1A<X]*;^OW<74 
@7TWU<P*YFZ!M\CQ]A#1 V5@ "P'#Y'%0TK$-A.NOD4T 
@5ZY"H+=LQ)C<D 5.G1_!MSA,<1QQ/80BEW$E$L"F/OL 
@TV84"$6\2XD):1]H*JY U.5!FZ]B'%CP*5/O(U][[(T 
@N]T^7>X6' J6CSZ^!__PB*06!CX>@* B4Q^&GJ?J_;( 
@8%_7U9KBT&.6!)+OC;NPC//D%@A$S@6.7[/C\(<K@Q< 
@/0JA-L>1ZZ/N\,K!]!R#T8P(ORLKT>B#^&WA<->";4@ 
@K^P[K2W$=?47W J:J:)"GL4(]XUU.,D%>1R24JWPC[< 
@I5^X&C7X52Y>#BFL<T$P#  V_\Q\?C9.R3>C<4_S0+4 
@3J'?7H5TTGB,AE2QF-%![L<^S:PB04,+"+QN\^HLWJD 
@V-=2RF&#O6D)FW@YPF?PDT)_MI>A%H$J39W+@8EY7'T 
@MI\<$PM;<^:U$XU<1N*]I&&Q=N8H@-@NH_W1XV:X!I$ 
@&YZAKS;<"+[,R\N<>2Z;VP,];AL)6Y Q3I83=!K;\!4 
@ZNW+<EE1)2?_ [_-#EV$))TN(NA0T8.$N#5M6(G1YR, 
@Z*H/<V5787+J,M!RLFZ\1$F-L,UJJ55:<1"%DDH5?G\ 
@>,'""W3<"C16VF>Q&W1RAI*P3&?RUB#U 7$"C0S.,)< 
@ED76U^]P#O3G_E\&%%?!:(6Q5G<$)G3FH8^Z0*#AXV$ 
@@IF MC?UL&1MOTRDB; XO@QW$AY<P/Y ),87'<(EXS$ 
@O'&P:W"MKB$0&C]S03+ EH@3=5Z16+Z =!_X;_TISWL 
@S>OE9+ZH <\^9>1AQS]; ADP='<L52Y)Q@&?O,=K?#T 
@F'$-77VSM?O/LK.-(4SJ]<JEVV!7'9>NX#A0<4=+MX, 
@A!.[-^ZOBF)7@TM!\2#F\\QBZ!P2^G:ZC<'&B0.^-4D 
@WKO%5>7Y)2DQ,5B"*K^X7XA4#<4=F+;'F0DDJEN3'ML 
@\&6?"X,BP71IVH-"46@T[E-URI26K&@&ZFZUI9?))VD 
@9(D! BO(7O$F&MM20\11XR*RSY=[VU4 ;\,WJP$-BA( 
@)3XC&0VFTABQ3OGOP^[==P>(7CE]JQTMN!Z'>AR>8>( 
@M)<+DAVP'6_*S% #WDF?S]V[IP.YN-V:.,N&7 SP*)T 
@XBV43]"K?G@5W6>\=E0+BV?K=,%,A'GMD2_C,;@/S%8 
@=5"WT@M-WX2"9SLB5"KNW3 K9)4&<QW#W/P\_SYKW(0 
@3MW8T&_X_=<.4>Z_55IG9BJ059Y?M;8G9M[]0]^%#6$ 
@\[>MH(ZC9&Y0_UZRN=?[6 L?9;L*Z2D'GSNK;XHM U8 
@7 &1!#C^RAL>S5D12@E,D;N#G&#C G,EO/XY_]=_S"D 
@Z&-H-(W4 <RH)26SX2,;XE$3CN4I,P/P#73=6/S4@_0 
@4Y&WA4Z</SK.*VG@\WL6D_F%& F(7*P6EVFZ3EH(OM$ 
@5M1S&VUX]Z%4265G &Q=@*U4$>V!%,)4D[V"BR%.Q,, 
@J"1D)KD1WU;HPREJA6)DR9XA[R; Y&K5WEP/LJ+^@[  
@!;H5NNUV)QN<OF5^W&XD%3H.GZA(-9U%K#%\)V6IGGL 
@=WWJC? 8&3LQ&-CJ31JD_!D.T ['UUXT]A3$3#;S/JL 
@*4M6:W\90Q&\@GOM(/9&4G2-U4QN; 0E]H6,W9TN^1\ 
@J&?8XHD@(2>"JQ#8@"6 C>1)?=OC"AEH 00N$!;961D 
@M!U&9)5V?.%A<R7-H7^N$W&'H&[H(50NB)KA3X3&>]H 
@K2UE(T&P*Q'^7\H':%@FTTN:!FO?>LIA&W=UU9A>!]0 
@+ -5./TRNZUYURJ#@5/[4OQ\NJLD+]?(]XS9WI&J9RX 
@/J3?<UG!;,841 %.;@])=?<JK0RZ!W6%F]O2YZ2+_Q< 
@<PVWYU:);[967'[&$3JR.\?8 <02\6X$> *J2WPACW$ 
@VR,SFQ!14 .;^QV3.\P>7#JX>QZF"IO>+KZ_>YYFLOD 
@%E=[1MD^Y1G])I44BDCO)&&A@_O)?O"O]6D.VLS')F( 
@83 ;K)N5N4T@>E!,';T",$'NYQQJM_.[+^W;#RZCP\8 
@HE[BCY"<L=#T?$>K/+,?*C-G1(C[/HWXN!!$G+DN&VX 
@>H,L<)MR.>'F+6=GH*]7HQ0Z&0P+M2=SZ*2/1] Q5,P 
@?D<AXEETCDU,5(O;';"SU^*M!:X&=-SL0;9F,7!$#(X 
@(1EN6,$B+2I5%Z"LAA#,?[> WQ(2J^(!@WL&D(NS^V< 
@#)@A:C. VU<Q+*$!/T@#V=^2#+R''C.]ICN]N\8%E8\ 
@XQ\92+COSMP*8HULF>U!5= 8"8%LP<\$BE?5 _K)1$@ 
@3FM>R)N82[K*'6G3:\G0=P7)^#((7'IU$@F*[UQK93, 
@!IC,P_J]104/E:+^W17FV&)1#!34;4_\'>3&T]\">:H 
@Y<:RXSJC,/U(3KFT!4">;&7Z9>C$7B\K$A4$MR?$1H@ 
@9B-)G/4:>U^M-&]]E'PB??3)-!0LKR,4ZW2,F ]*#A4 
@!=>"][GK,G#O3%@UB?[LH2YP#]2%Q<E3"ELU_%&S:^, 
@[J'SP-?XG@Y)P?G\L+=C@:IG1[:.>[.TJ04YVDP@NS\ 
@@'1E"FP]ECPRB<HT&1E(G@3+A%]UM/(#^=W6^5BZ*"  
@? B!S-&M2"3<#VUP&+F^RX]GO '&L'M=?QIK $ 6%4$ 
@2\Z+BH'IZB1BZ-=14R5D\[#9KAE6[T42QM6N=NL%8E( 
@.'>TUNIIG]86K1*EO\RH2]_8>.<9 &C(3T #H!,N3N$ 
@WH"V5 -N\_*OR=)APD?\5P:#Y$]TZ6<[VEG\SMM6+_0 
@.YS.#<Z%]] ?Y"DID 3)*>)#W87"D.<TB0H,C'&HE@  
@,7!A'1O)@DNQ@WXV#_LX>;O,4)$PWP2J,\</K;UW[(0 
@\^6:3L^C$GWM)"ZX/'BC2YZ7<XWRGC!.]DX?U?98+I( 
@KD?@BW.!]]I"15+73^UE*N! C)/%\4#$>4@8QA+P9UL 
@A"_KU,0C"5WRC(&WI;2ZR^7*]R: Y$?RA(\2&3."[!X 
@@U2#87]P+4-XB[G*;(XIP7-OF(WUKB4!KPG'R.@2.<4 
@V'FEO<V;.2T0#8.VUHP!JX!/KZR!I&QW;.EI%EM)+(0 
@7_^%84"W\_W^X)@F\-%E!L>5,/Z*IR*MAL?W'YRT7]L 
@@F3:JX]$G,Z$@.#2G.-C&C!? ( L15',O#9#D7.J0(@ 
@: M.4Z(8H3P\-DSX? MDS0Q/5R%C)X+CYZUW]E)@XVP 
@8Q+D6\AX8O&LP=?I]-A))OZ(HX@XJFB_)CH3K27GN;$ 
@U;=/$$/A2]KNI%H&['<B,//_(?D*/Y$#\/')<+=:124 
@ZY7Y1"4+*YWIK;#(TG*LLQ_52R3%(E!E%UX<+L>MJ-X 
@)E089TC/JP.LIX2U9V$I#M%?QOGK;EY@#9KCXA[CL&( 
@I\11'54AE2$2[0B16MT0[XP.O%ZKH91^3UJ1,A8^",  
@>FDFBU<()1CSGT"#01DQ97E #UGTD?*'U)V%&'JM#A< 
@,N#)U_^1:=T=<)-9U+2ZW7J5_!&!@!OLS.KS.U]RZET 
@% +7_XW8;0MA]>FM[MGI/VHM[:J6']%0#VA'2BO_>(, 
@X9A5!25_W6RW6G'ZO*FRN5P/VYOQY,Z>$2QX2JX0#;$ 
@_%=4!Z?0N1DB%0.)?TR%LYR1V@0!HY'C5!K@\<$]4.L 
@2!XD7(YA^JLR%QWG1E\5B@(D=3'2T;KX2JP<R/#"B2\ 
@IAB[GUN&3=!H-.IXYTLQ2U9+HCGN%10K>8H)9?CD$!H 
@DDY[=P[%>(TQK+5$<>DF_XFZ8%_EH_Q-+B)^55N<W1, 
@;>ZX2]O4>M.XQ.2-]=]402MJ]\AFV[1N%RW^'<>D;J( 
@O8X!,_%=!I/:?[+PD]_TM X?&0RYS">5]H2T2C7H4<P 
@O56KA[@M313>AN4>67O9P+R=>$?=&Y6VK+ N2UOO*3  
@1PK'2ZUK_0A!7]*_KL,MR\*O0:KIRN"P<]H4C_ZVM[@ 
@9?#0>[.OK8*27PYZ42-8-)! 2.5FUW+A%@MIA7W=ZW4 
@U6H9IQ\PQ4<$B=K#B&@=NYJQ;N>ZU2EY,(-X^"BM=>$ 
@]V\5(OXB]QK(V7TK5]8V3&DF0+C9I?#F -J=8&UUIBX 
@::0?2=U+$WQ'^5IZ4X9U],01,2K#5+#X#JU- W0:(H$ 
@T\YS"](@GK'M&!.NW+7U$Z$KN:7&.LI9T$NJ6$*JRY0 
@R*IQO)>??^8T]!A9)RQ!O",+M]*@ 6XK=WYYSTM=ROL 
@IS3+0:[>A/-/5<VTO$[NVWR; @!C@3*O]_4:W1T[]K0 
@. 0<BNL"%4O<KP.$QJ%O6N8N@788:N!"E"8QHQX ),\ 
@?'I[XL877D ?A'/[IE\PM$C5V]+KN'V83"8U+',=(;D 
@L8J_M$5\A*_]RA/"%_!*F)H,+U9^QY.TIU]K:-IYEK0 
@F:_2(EV=A^@QY\D^M6TDZ_8GH: LOCY3*M^0P2Z10YX 
@FWGNEH._SEW>Y/0GW32X23PW##X5$^<!9REEBSYZ15@ 
@]E-WG&R !TEW1SA0"H=#?*@F);@[#:G:-VA,+5KPM%L 
@M^#X1#W+30GRGZS&4'<M7XFX!WG4P<PLI5I7^;62TD@ 
@5-/3&Y?ZFS>M:3:X'?<]']G+"RFCX09I7_'WL][+XO4 
@QRE]00;F/Q@K.%W'M(-@@55Z]X((QCS['+>TMA)>%N0 
@X .P4,U1Z.D9[&2ZD_XBWSB-%3AC%TERVF[]>5I\[_L 
@EV'O1%#E )W-K%GA:&J,!-+>\B9MU/\CF[$N,Z@1DN@ 
@"<%QV%-C*TR#S:IN-E'(4Y*!UR>=]<\>XJKM#+;R+0( 
@0=.DQACEB7RO2<>8'8I@EN@P<N:UTK#(EOLM1H4^/R0 
@+W4D).*]R7WG'< Y?MT\9-H\LE09C(@'(W%+P.\4_SH 
@]]W_4<SCOKNDCE.".Y,MD=RU[<FA:FM.D";JB]RD3-8 
@&TNCDC%7EBB9:PEAVVA<H>/X:+X$T%@)PB# $SES3,X 
@Z@WTMY=H\!#*Y$6X>1..T4#(BI (.9=L/!)?F?'MCPX 
@_NKUQS51<#4>L5O[5ZEKK.)2Y?5WY;L8_X3O.F4X-U, 
@0.C!;E@VK33R6[R1#6626VCD#=]LSKL856CERM*\/[  
@%MKX)_#78^?9#B\ZQ TW=(1?M(0ZRAU$\U<^P?Z\'#, 
@D/[K$-X"[*')/KL8HM 7X(0N.B^BBRG$!7L=84ASAN0 
@;C"%=PI$ST/A##A]CA)ND:W]C5+P]SV2U%CD96(UDL  
@_J 2A+;;08\D2*#B7U2W=J& 9-JE3!^":;IO3&58S4L 
@E8<EADAR>RF0M>\OWEXB=OO9,$[J0T298)6JC& HMED 
@'T9*OA9[U/+<QL2,=](P&$K:TKGMU>8JNPW]MD/IAF$ 
@;Y[C^%,\WSIP2GQWT!A&[V(@XJNI>&35"G@U8XE=7[( 
@FYU$++5E#S@]066,+G06171OPXRLWN1WF.!G7M&JEI, 
@YPSR8E6GHR4$UILN42:9+Q[/LAH2F5\-.:X4JYZ>+_\ 
@F4!CR50@*:@IG?Q+RH?H'C0V (UEL<[MW0WKM8\]7WX 
@K_5T(:'D\QH%NZ[)F="4;F5J/CV*VF=W#D!!N$'R?F0 
@H^LNZ/.K![V UT"D60(";^L=6PVVHFGR:F6#5/4VE/P 
@3L/O)WS%PAB_;D4'J]$LV0])'R&)^1PA$HYK5M]MF\< 
@/'K.RJ"%3I>\DY4HB*GI@FS>_;&]C\+P<E0_YUG01'T 
@>RQ!/"Y5A0C9KC,F^:;^)K3LMDWO(<6E127T![A=0Q0 
@D$5O3:>Q&S:7%;!KK@:;@H_[?* B1;OA\OUW'MW5]BP 
@QO<JECY)/8F'8Q8B]@M A1@&BU<4[-,P(RY O]W?^+, 
@KGKY^)/ !&%KAJ!<?\D7'=%6M"=[Y,S.[(:1&0GQE#4 
@8TKD1#B:)MN/PZ3791L@UI5YN?C7%1J/AEW/S=:?SN  
@G,QGF*ZC>EBXN):8>*SU7- 3Z6KY)E\(Z:GEI%5MF^D 
@V3FXW2*V=_:=Z50Z9K+)?[F*9F58CF[8?+"2W38L*Y0 
@/*D @7DT5TU9MF.LOSY!MY8=!AC]O:(_%]8J0Y*0])T 
@4U*M1:%@WCJ""/;(BL&TW\'"0&'AY2!B"63Y0DAFYO8 
@>1<DADW$8E*KE79V R_C'#:?6I=LU'J9MH19N*/(+BT 
@A!,A7QT.YH]XW4:>&1$$#"O9"C_*10? N:Q+"#\_+QX 
@T5BLN,,[7L-U)2?DV+Q@&A%1,Q,>"QJ:;(P*)[T$D:( 
@PH<=+G14P4VB5&S. "2E<E5ZB*LHU5/T$X*'W'QA?+P 
@;W%BSDT.Y6T&RR$&2ZDZX .MX[?7P(1QB.Z[G:@#\$@ 
@WYOM,B_"LRK6/L))&ASOA+G[;T^#_37)MKE8V_QSTUD 
@\D/#P.DH<LYX>(:+B\L(Z<8B!"]S*_;W<JR+T(_^M T 
@VNKOO:PS^%_4\.\18X&N+0MYP&>/')/3HK:SM#3'7*8 
@;1&%;&NN ';[/\'NVPVSDC'UT"SU<3WL).6B,W\A&)$ 
@E!@$4%ZRHZ0-K:@@Z9D  U+4>N0O:!0,B-8V2S5<_CT 
@Q:QG ?V]]WV@/EYE*86M?FZ!ZUVRS>M>-I1A9%.TM8\ 
@WQ,\;Q-51!BN<7B'K\,XKR+F[$>*<E$I*.%8NI"*+;$ 
@>140!4B82O)(]C&-]0V*]=O.6P*XNH4\3(-[C:MGH)D 
@0G ]Q2B]XP)0X*;%>N7:&)4&QWXW"B<"17!1TPIIBH  
@:-CCIE7S/FQMUP7#D!&O3)-^;:-NBD4W9Z^5+#[,6!0 
@)N7[4")"4+!-G2 +^_'7J'LT<6!5 (*>,S:BD6*3<8< 
@IX$L",^CV:=H9WK_ZB\LE%:TQ&J"MA!*2T8<4)/^1:\ 
@,[/N3OQIMR"A<)M__-=<K#,9/V\BNN'_IWZQ#5[62T0 
@%NJ1=FQ1N?)[,Z="%$T"G)@SR^,G"&!'TPY+A^QZ<AH 
@:CV6"R"#-L&' WP9K_0)1_I0WS90BMO0OO:K.\5X>7$ 
@WG@X(R?$QH:4NHIXOMNF7?*;F4->3#=V!J$T':UM=O8 
@>(FB>(.M_L;R4F\+D!T/#>,=\&KYUS5>]"\45L; 1SX 
@NOF%JZ\Y3ZN0A<+86'IK54@O+;+"YA>_>2>(+_S"V^< 
@&<!+&]G_I:*VY-G/[%50"-&@8>D&;>R0=K !681@<"D 
@J)Y2:8UYU2VL>UI08=.,3Y+J[O0__J0Q"6?_5]Y=2Y  
@BEU@$OA2;A4CA<65+:TDNJFKG-=6%!61\BV5(;G(7+8 
@I-!^*I0D=^A4^D6NKQ FTW\I>[\VV5.\%-Q0TH,PF$< 
@PWLQ/Q0W@ 45V93;U!0SZ8X;J:.9<$^-I7QQ]TY4K7$ 
@W4EZ8V7&C+_!)?'HTYB-M<P"5URFW <>H4_"FJE9$!8 
@6!$%>J$>H7XKH9FG#3U"X0&.@]=/BU>%6)-$_<"17'8 
@J5X\MC*'HT!![67VH+X !2,!ZS7([G4"=&\V2F^>.^P 
@%Z?BL;S-!5.8[@+8F9+B/"\>6A:D_T(6'G:S$D>@(]4 
@Q4NI9C.Y!OOD"#]8D (D;. M&=ZRG/YM^/06]FGL#\\ 
@RT.0$ZIE,+ ]?-OR9C)* OYWVZZ$O'$N]>:*PG8U:A, 
@XS@CZ\)WG&9R/!@L:.;&6;M$^603"Z*)*_)DXP3P!Z@ 
@3I'_YL[T)CR3^F5  (VX:4?KL_G^OS.>OHT:+E[[,*, 
@JX.$-Q E$__>E>N+V7NT"!.=OEF4^7XS9>9'$R-:@IT 
@_N758]YO0.LM/0W#*S]C,<.QL#Z4E*/C0PU(;!<DRG  
@FCC*X^7R,P @M2GMRA><.6'3.C\?)^Y]%(#)C9Z1#WD 
@!6.1CB\@&5NT97Q-5 E.C:T">1'>\IF$^-]&JT1661@ 
@CS>!A$/LGJUEYUWKLRJ%1<0%C29M@#;S0"[+6HIE=2$ 
@E?<0,1R S&- 4?;L-7U.)A/4"I=7NT/Q@C<G/FDJP84 
@])A.#,B:Z(ML^^)5&A!V.E*NG4D@M&+%OY2>BB]X@64 
@HNR&Z2+ _D9V)$?Z_'U*NW,_0_?UAKEBW#@[) ;IC%T 
@)5!'"WE(+>0,RCFY'@YQND_(2&M3.\RG9$4_:34INOP 
@=TZXFJ8-<.VHG SH8O]K-?T:7C*DE<,<K[N<O[@Y/?H 
@M6KZLN*J70.N!0&$*TS8#H*O/Y!OKPVN3FV.CTGGSP0 
@2?]R_K[&1%^/AP*:CBJ[X0\M*#15JJ-C%*H>M]T!COX 
@#S*#V:=0GT3%VY5=YVHHKYX,JXHT&(SWH<AR<?GLHM, 
@CZKS=8!<4-S^EFV[R?J18\-8NO?PUQ=$X.6NC_^X?F, 
@.C6:EF(O*7\ &.3H/EH;,2I157< Q7/'DS 1?=&JO"T 
@1^F=O[IEH'P[_(T0]JXH?MCU?8IKMHV84KG("!!X+JL 
@@#V%+CG=Y5+6IK-)RN\R@DI;CHQ&<^";.W/,JL84. 0 
@(,?@Z&AD[YG9\XQ#GNG?O^XTZX!VQ4NS ><=#8J!$0< 
@3[PP:?3]'Z;?<#X*_8=<P^@_J:$Y2[L: 6U$80N*3W  
@)<K/#F@J)M[L$2;5M^'M9)=?[4ZOM["'\ )D.#W+1SL 
@[J^V?_.BJ@[2YZ0Z^  L[ H@NN^6GZ,Y=.G7>8==6DT 
@O*.*<_&Y=7NYCO^DD[ZTB#8 FS&1P\'M+"EIGTR,"G4 
@(#FX-NS]4$\_']NCH?1GT*P<I>BGP&GIFT;96*%E;-H 
@>$NX45N8OR-LPB[Q9&>.JRM4.4UVK>1!B' (CX79X0X 
@NZQ/K7K$]<P/#H,0>0C3"$&(SH0W60R6[8O]'MJR_:$ 
@ J%3)/! T*TP-C!E^%OWI7A#&VX.!-61L9?F9DO2.CP 
@Q.6K1\@S#=FXHCB-[M],J#YLF/<"?$L26U?^!L="RF$ 
@V $_;I%UKNKBS,FD:K9<P#3"(..%*2*M2V%K!K0+>4  
@CBFO(DV-S)/X:;;Z3.8$9?-9W./ D@J.]?*PK-)/<G, 
@[>]*9:^%/_8CK\9@6L2KJN(&A.X+N];#MDXC4+Y.%N4 
@5?.G9J<NH<X%_7.O2K\<[P? M%')P7"7L8 2A-VTD,8 
@)LSZ?R6;VKN8P'\!U>RE<9$GC%KE"?I)'EV\E7O2:*X 
@N66P'[9O@]; 5*!F>%Q,[N/5H +%5BU'4_*O6#^VY5< 
@.IU'?<>JT-@_N3%)67!$8Y>^>)/?5_Z_E_V]C@8U4?, 
@.J#6>34Z<9EI$,IFQ=0-_+;55/M!M8 %2B&AA(HH*1@ 
@G&+-<O$G\(WGH#+ Z"M%0 JF4B68C 2/:#185E(ZO28 
@:Z>;!$_(,YE(,C<Q=CCB =_LGBXU-[.1[:@CL] F,\$ 
@XP'S:=.1R!;/?;UK-<J-2VK;CM,O$"/F-V25;Q%,;'4 
@?OG7:-A>NLZ^&<7YA,_BS01%!1IL8$O,3HU;0&0FBO( 
@I6:&24E\WRXCI%]$FO)KVAJ$L0MJVV@D P0,)GOR0[\ 
@'[ST]3I(D1I\CCG[1;YJM>SLJU!<J'9YYFWZC1M/J/8 
@^)%"Q2IXB/3#B?W%&.O&=GWK]IWV$*YL 99$9R*R5&< 
@%X@/D)*UUFGX:0&-X-M,PFFN'B9.[SY",,1N.#F3?H  
@3I>:;. _;MA]SK$$:H=OA?7BXQ-<+N_Y$H%L9*=ITZ( 
@1C;Z+$7D^]J@W7=NYG*KB!^NY>#8/C"@.X\DNE9CU_T 
@*J!$7J2=MUOX71/+=\!IF;5()P#[V"A,#?/^)P-OS\< 
@"N@0'=,!R%/=*?38Y<[]96]PM]2T=S]%)NI#3=(.FWX 
@L\X7!ZL0716G>O1,+#DO^PP5]NRFVHIX1[Q:V03MD5L 
@'9G_['%%0/9=8%L)&L.Y/Z=U19/O[7S0N>W/(J!Y5*( 
@U<.FP^A_WY+.LV--*!5%:9ZT';]IPM2R[LQ%P&;#K&X 
@G/.Q;A6Q9JE=SVD"DA@>&2X.\L,(E?J)]>QG:[P_"I4 
@+<P9#=^3C/9I#S'];/(X^S/LRN<SPQ1(F9X4Z]8XOF, 
@5? M3B6V%T[N#T9^<%!/KL,I&54U/[^.%3*7A73>]S@ 
@;B]M<LW>2[H+*$Q, U7#DSR-,^''SUV?[Z38B'\7W<4 
@$N>(,"=Z#,.'OFX%-T/BBEN,+Z+4<V0:Y/.H@NL]^-@ 
@6HI-)_ZFOLBY&)SP 322/JTY0)*[A(PQI/GIUL* U@4 
@CD>C!78F&[-*7YC2&5WB>@,;=SY<(?-)R)NWG$( 'L( 
@=Z5X_Y?]BF_^\X+3A]"..\6<QUR;^D#;"7YT@YZS6(@ 
@?V5]$?P<93XI1=N@:2L[)503<<H49%D2*RYNI/<;P"  
@#/3.U^I>.AX:UC9V6*+UKF8)I&9736J1T*0.!. :[8L 
@H!HQ=#+R;L)P=2B]K0(BX99I9<"FF1>?AVIS2+^B9+\ 
@8DE9X2RCO0>68=6DF2Z@,E8GY60-<?C:' .I_OQZ^NP 
@1NU2J@WNH=3P-#@&1QMOL6I?"H4/N0V"HU?GJ=)-2ET 
@@;9PPKT:1MEL-$@.*.FP!8>PY=1&4]7[;]%4+F,\5?D 
@,\.7+#%8J6D8;S:#CU85#+):U188F=@5^4E".C$EQB8 
@R,1ZO4]_3-A12(:7XV^H][E058SY3 X<<OI<@XO>36$ 
@<@GXW;OE!&EA@XC[__/T(8.:@<AWV0$!;PJQ"%HMQ9D 
@HV?-3'^A/@ >N4<-_-7F88O6=EF(-]QP/:?CPGVTTF, 
@*Y_=C0P,8=F["/S55*L\7/&XGW?KRIC%:P&23/9AN)< 
@0F%:PVPV+2<,J:LT@LS1[SW7V7!0VLZW##)0NZ+8L(H 
@JVP3<&:,/=B0&D0%TQB"Q3816H]\=*>WOD,IBUK'DSP 
@?.">TO7$LH\#@#IP>7JH/%M,M,?/78T@*96:3CS+:*\ 
@!!8J?C"V92M#= #[31/!Z-":;L><YSY !4</>UMGW"8 
@3S_%9AN9:]2SN (=&:I5"-IJ*K&,G_:OE4)?RPC!ELP 
@E9>!K2*8MIGO]7"YT+98,5!;L00CV- S-HW2U#G_7!@ 
@M/PW.Q;1B*2;.OG(96V.C2-F?OB-:8_MA;0\Z^,KNEH 
@4J!T#-;[8)D*HC]^\?L\:'AP"_0UO.$B QJ:?2RQ1., 
@;/72:N+LRB?THK+V-U:;/TU.JK4RW%""F6M9H/CH4>L 
@,#TW3MYCD/(VXH$ (U62BC7:"IGPK05P,YMM.#5!+QP 
@A1F@IQ.C$H":YJ4$<.[X/3XCE/AG-5%,AX?WNMPS'#T 
@L#1&\M O1*WR5*Q7AJ[UT;>+GS\P11\62\H.YS%(1X( 
@;$C"#/0Q:515&B$/Y4%6,)ZM**9-)#WXRZ& 7P$(S\4 
@U(YF7_3YHDCT:^ VTZ-@="PAWH_%OP);HWUCSL=@!ZL 
@PNK3/5.Y/GHH/J;AG1=PQFFC=6E!B,7H.+:@J>:<A\8 
@7P8R#5(U_G E-*\#70"U*3W]*,[&H$3'L0K&2'H6W*P 
@9@-GU50_CM(W[]$**'B-=NRY-!%ANUF%BSKW]LQ[$^$ 
@?6F7I9U3%$&#CM*1ALMRA</-.!#?! 2Y'<RUSV1H7YP 
@U."JY^22OZ=S '4ER=F'%57D*E*":C"0IR=%XC]CK\\ 
@H^P\;"O<0_D%D]DC,C9\&)\E9GWJ[V E1CER,SE>V6L 
@*!Q\Z9FG'*?%$YXQ&XZEYF33Z*L5//@403FQ8SL4#U8 
@-1)$>KL_=@"?@EB+^.Y,%Z]ERZ:^3@*2&#5]3NBPD^X 
@:SX"2&=OG=!Y.RF4<U*\/SU1FM\".,DS$3OU9!%:OLL 
@7W>XD< 4)1IA?1=@L"$W/2P"0AKS?84)]B34+MYOR$D 
@M33-\PX#Q7T:,4\A2\=\0]F(RA>(R_HA%"GL@_MLUY\ 
@R5B"&6I]&A39!>*+((L&[SCLV[M;5]BS@CZ&@V$=M0D 
@7&SN\&]#4][KQ2V2>3B1"@FR/8OF%*M5X%M@]2LROUT 
@]GO8REV0?.K_E3*UU^$AU2 @90TRD,WZ*!TY+YKEK6L 
@+3VC(P!&;HM4;RW_0W(WYT&CYZ5H:4[?9;.P!,T8@Q( 
@;)=-=V;JV)!@:]!1IH;\+\XD5UQZ#"9_;9IY*GEV]C8 
@@(D4!S2JN)%N;$H1-D+M1"$J2%.*W_&;0X=FSK(CF>T 
@/F[+NR^S$\SA5*D!H9K76<OCZNO+M%I%)'SH$WBU7X0 
@QGLZ>F3U=LJ@XS)_LX4$:#^T9QN#PA5' = D!DO)(8, 
@:=7823,W_GK?K05/Q<@.->^_4!)-.NXBJ1L,_EXW-4  
@*"AV?1/?<95<_//YII:L^9).''TBW%*#*%Z#?;4?J9H 
@=A_P]O^B93!D3D@=. U)?M8,M+E1<Q2S4N:RI)^80-0 
@?4#47)X0IEI^TGHDZJ9.-<I>$C\*JT' D>!*8E#(34P 
@1HP._EQ$+GT+P)&NYA&0_WQ"<^"$9?[&.?76 +M6NQ( 
@Y]]9[ VX5) /4733',W  =HMAG_Z3(NZ:R!O=*!?_:0 
@K7\]U>(S4C[U5EZQ25OY.@QA*9)_%S':483R9[]JUV@ 
@P#V@3*ADP>34)/^1B]\"7E>0$RP4O<'Q55JHN0YBK84 
@SY9CFE['W%7Z:2PD)4LB_&655,O+!&4&6!XR*N?(_A\ 
@1"P?#.^O[PXYJW4 A<[ZLD#_U#L  TY'DY&'DT=MHZ$ 
@E'KM\ +(P^\WC)?)V";C>4&)8$^.N3##3C*8M!2.H?$ 
@GMFJ#NZLPFCWV=VMX7V]V4C* %QN%(=@J(2^G1 L@DP 
@--EOB,-ROKYE>':O%VYTU.%Y*OYUY&SC(M"-*YK PVT 
@;_J^KK\7H,?9<&=XL]P/7P'1]^[SJC;B/U@5[U"L:.< 
@TQ+5Y/8'E[X]1)SFSFF3CQ>'-15XBP\F*(/-0P;B:NT 
@U0$$A#3YBZ3WBNI=HTRI'DH5X6UDY4][L:?:NK-A'^D 
@A+AU-Q\*G;VD4D7D(NR\EF!7-D@22_-9<UU2\,C8D0$ 
@_"B_2V_^\%&_6^+%[TU[2!TNR06I6QCJBP!#"C03^0T 
@&X*54EPD>\(C^R"S=1O'M 37ZE@X<4PVE1+5RL!N';P 
@IOGOYM!<MRF$4)Y^]@:Z DYIFRLS,@8O9>7IQT]Z;]( 
@7+CC,HA7K[L4@*#"XQ\(-]?%E(\8'K!GY41JY*$X1O$ 
@"UBO?$EQPI_0?6UWCN0THE^I^I/M=[PXU'O)(*PW6.H 
@9_C<T0)LOK:2"E3FM8+T7?=!%R%Y",RN'I484WEE!L@ 
@4SN(4L\C<J"B&Y9C@6LLA$4:U-,'=]QR^ DRWJZ19Z4 
@('CQM>X\AX,\<0+)!MW7GF:U)BDD/R?9$2D!N&)Q$W, 
@=B@JQN?KJ7 .6&^ !1>3SG.&+;BY3/C,-/Q!R"1B='( 
@$H?PWXYX'89P]MW7:K1O=JWP0RL#CH4.T9%<X1C-%40 
@:[*<^^\]D:)!;Z1)Y\_"B]&(=K&LU_P$<JZZ5( (*)( 
@+ZL%2?>^IRF=QAB^J)>?<$S?:)BE5A#DMMFFMB@:?;L 
@KKUQ&378+H!BF;S#T#X@9P Q<+&F_9G ] CPCY&E8X< 
@>Q!W)EA.+_7>V(*FSR>=6IVYCO0L?,;:X&+?"(1MV!4 
@*W^F(HR^6O<QHA.H[D<9TZ)+HS6=0A;MJ_#=Q425=$H 
@2ZDT^0'-T3A)2$:R47TLD+?[(T2Y@1'57N'P>8T25"D 
@#'&/NM,.Z\6K-6U<)YO[+!5:279G*2]/J\>3C%6I,%8 
@E8\:0G:"V7][D03,-QQLCE^O*+"0+W+XN+LA,PQ.B'H 
@\FI'N80J,=.,I ?D@P.ZQQ-8_&B<K/@A&2U=XLH$114 
@G>?VDS91^AH9'-1]O ]5H([$PIS7?':X;9;)A38NT6L 
@^>8^L^GY<K;M=6VLBR)).P!;7OO:2">3&[I%0KQ!A-  
@N/36&?F-=FHO8!,E=%G*@%B.9VR,V%X_&"F(]^;,W8P 
@5:F",D<S>.LT'GIVIKLN9#ZIRW-;#0;<I=.E+1"S<M$ 
@>=XU!_^@LLSJX*R5^H[1Z#Y\VT0&NO$2!#@;^=9982( 
@E0@G"2[[Q?W22[#B:S$@G;[%+.HR&#3(NB"D 2] OOH 
@^ILA\'\?"3#>9N!]4N>":8FG<'F.\9 @[>*^76L#?XX 
@,=/Z"P_OT@Y3<\:_04Q^:.>+=V\=FDZGUT1H-6E7^!  
@? 1U38QI.LC4WNXLC%/($+BRD4$'A[C"O9\["G\=[M( 
@%X93/E]MF#=[VG,ZR62$GEG(J'_P.]G _. B/*+L0]4 
@_.+6'JM>T,+H\: 7T(_3>48#/5Y"?NYG&?O6$:KSI<$ 
@"73RIA(>R$!RN/-^;5%2*"*P8-^15V2IGGMV/IM01TH 
@6/W7N]HG30^DU :6>G%22HKA:(/HT5M?EBHFT)!-WO\ 
@F(@:S'])64H5H)+XYP"'"@C.!!.RI0.\3: E=E%+\9H 
@#HO?0?4HU=A?R"1"9A$_P',;V1.62+PEK/K%^6^[ZHL 
@S?[7YUT,[TNL(7JFZX,^$,GN),D&&6RM=GR'U[;<6., 
@A$61/[;%8 +NGO*:G9+)3G.M%5L EB!\>FV!&EH&:5  
@C QK :&*SZ*3=W?T=IN0E;)/T]0IS*ID#^Y$UP(6);X 
@E?0<#:N-2JI7H:5&(_)O^G7#9T," J5EQ>T1I#A-1%( 
@\";58Q*T?JU/?%F-KF5^SX/X2M:47_?U-+AA%6:8VW4 
@5^D=*9K#OWB<Q[2GXH<*VR]5^$LKH(,$8[6-Z]:%]3< 
@7:QJB<-T.H[3H)S6][$FO5)ZO3$ZH4?VJ!SMY)DCTGH 
@$R7M$>;39R5Q0X_YO]+GEB+-&3:Z36S)7;Z6-FA[PU$ 
@TSA%1M/^NVW)1QC2R[\L5)>8G$US[O^M*&$TG;'NBGP 
@PKB/Z0EG?.;U:I"R#B9?OF0&?(V(?<!1,;TR=P:W/@T 
@%!J]J8_<XC0$ LV(]%N-KI877P8HV3ESG,9*TEG+TJ, 
@\[FG:#70,?"G%;H[*P<[4/A'8-CB'^L?:_V@[<(A0XP 
@ B.*):3#1\@AI12=:8"/Q3N[V$=J5L\+VH3M,>H.^9( 
@B#D@DK?YSH8;K&2LMOX4*]FSF<2II->R?/6@V94[P$( 
@N&[A1:,7_]:&Z&P(D)%/?-HB=4:]-*'0DN:U\7@[2($ 
@KPUPUJ8<15'4WS;+Y#98% BF> (SKP=6LB[)=T,!".$ 
@OL)K9!$D]+7T)#/_9ZR+4N8UJC[H!,G^G.V:75/$KUX 
@ZLW@-5(K;W,?=U2[$S@KJ6>(!/3"/7/&=.PHJ[! B+L 
@C+S86">+ W))7U)+/&WSL/ST41JC,O I.O;M==[/84( 
@-K_L3EXA;./MH^6H8O(0(NH+I+H(@>+T1C&L5'?2\J\ 
@R$XX7Q49LY9?4!+^"< SCZ6JW2D]O=]MS]$?8&A54ZH 
@ F)VC8>;6<\S#UNN<^4B>/W965#;4#I66P$RB@Z7>;D 
@N%(M\*M1.I===??+?]P^$V_MA.\K9?TSL(\)U#\,I>$ 
@]7J36\(ON.7PPB1'2IE!^*B+5BKUO";_DCXM*VRE+C$ 
@%E V#=MP'SUHRZHY]3IIQB'CO:?K7( !.;5U 2)9R^T 
@NYU.:,"T_&\(TX6LKO[ \]WQY 5_\=:BZ"ELVJ#;VY4 
@@YH^%5JG_J>)+D8;-&E'>BP:%/0[&9H]N7XO? UFZ&D 
@"WI8TS@0J:GI(!,'=P7'53<=[I98EYG(3I)@O%$%!Q@ 
@VA(EX(L3P]\0CJN/?,OCPJ:I7YINC^;!RT&V0/Z@4!D 
@1#F7)XT57@OR@Q97HA,]H9BUQU*X$"=?(S570]H-3]X 
@ZUVYKLYIC9^[;C,)'D)F"4G+<P2QJYE>2WF^K8\RU5$ 
@#D)-8"3!#[3E!9_4(EF'T?\S_V"UV3MZ><0_-#06QC  
@VFXX?$"\)1HV]V!#_^!=B4R>^V]),C9N/3Z@<,KZ Z( 
@U_&*\ ^<<M_O27\]+5.,B<E'_/KX4+O8HU;]J4+$*3  
@<*<#\P4HT#6)S29Q^JRN3L0M5AHM?+=_.6\;B!5QZA, 
@LMO@UW :O*"-=GK(J 8VN._:*V0/).B'"W,"%^/I;5D 
@H<XM# 8ELV^YL3*HG]P>+[AF_L;3+X=6X(5%U?^:ZN8 
@=Y'!$^,<<]:?W$>;*T&B2G+TPY+)/?EWY3$%5]4?QF\ 
@0[^@ F.IT,U2^^[T?V)+TTVIWI>4,^KHQTS[_[DIWU4 
@X)1&X#8^T3I:(_&"L5_8? JUN$-A-;%YFUJY.%>X3R  
@'S\"U7Y_*<Q$*!7PQ'E-K)Y'7..?-FAJR\2*1K),%\X 
@N'':,R\W-^L#4,A>G7^J#E0]\$P()-PQRJ3\B>ED(O  
@V4X+-(K,X-=L8SIC&-=<5'1XU#?6YYBCJ.B!3S]#+V0 
0YQ#,3/+*&$X+1$^'F6=OA@  
`pragma protect end_protected
