// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:52 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
OOajr4nabk2yygyABVvT1fY/HvysPwmGZxU4i+ZkNWQXbrzTuJ515gxw2oUj0HiG
XGV3bS9B/Mslvu/Ka2qQQ1txGy0ZuvUzYT8A8kftpFKnHIDYQ4t2wyUCfcG4bKFh
IrNaRCe856z/f9DyQfLANhoKuzg2H7/b4Figg5ePia4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6352)
Ht/QBjafxFEag+eFh/Bl2XuMbaGrdaSGnjFLarlAhb2KduiK/YyCJ5ZhGOHDV/Tl
/lR3M50orDilIGo8ePqKRx97oTf8lyF1eMDVtaBy14Fqe8VflpNkhj9tuxQ0vqe4
R7AXR+lNgXwei7gOn33BS9Z/In1nxjWLGtYXCClci40mKLIXa9ATGQScBVXtdtR1
nIdPUHp9Lsxqm5Qga9dvyzTjKbHUYdpwfxP5UAh5S7RwjiaTEY0GaAVfjABer8RT
0oy9E2d5lGqE2fiVHDeTCZV6UR2aVzcPadBeXG18dCOP2k12sxN5lyhRwsfhzSHf
GQy0hO7CRjhXqGVHeMD9qdNYzcQStjliT4FcoxRxKsJRTAeVa0/wz3dMtm/+QBKa
H4TOniETBDHKTMa3S9EQFny4tO5+vzQN6PF7bRTYf9lDdKfvyMcW2vmU0/h4oMm8
ek4+6Ek3Xz4HRVPf0t1nLKJ0l9UUHT9SquIgOFRAYmPRRSJCBsSSEZc7Gn03XB43
r4ZkuGvK5jrZOngS6lOoRlavDB+An6w03ssbyx0y/HQpVZdGpT21hyE2eXHbu6Xu
vWK/jCp0lXF68TS+7h8cG1HVIcwE9Vcdhlim5ri5eAU/u9fB+2uyMXsPAQkjOVnM
hzfLR/orL1ufSjlTRKl72I3NzkgQ8CagExTc0SXbVQ2G4+75XW33pYrSKRa11Z+q
a+iUV4jqeXKTvpIiyjec1VO9aM9Dc/DUghNzM3oHQYfFS6aGNVFHMoxkkoE3v5Eo
D/+S4jvFN8PsVEdEAFyDi9o2ikmF3OrYqVp/APtI0ut+/oyAYhYaeKxJvYKa99gD
V1Bmw8mgkaHOfYjjHMbPghNEVl/85cdVWXgXxK8OgOCyr8mO8MkeGqi+ksm5/cUK
cdh1BfuBQzmIXfj4bT0UV9htrZZxJbJJYG43qNVLwa/3WU9paovWz+YOcjFVPKAA
iHp2PYYs5O2DRYmSBadTz/43jXusgzF1p//MksLePA2Bt8xXKJCfsEAfUFWfQ+W9
Cgr4QRJwotLa3wPjXmosW4JeqamDeBdeUa0whI8KRkaYD1AueFAQ0NYD06KrkUrf
XsRWls9L4sLJ0FwDL/BtcuSZElqUDaiM3Xp3NCXCenI+ZntHwq8b/Yf+F7Id+0lb
DWZAJzRQ3li35frOftsgY7/A1sb48/dS+c9S+0PxnYbVKltrARpj8PuBzHQVWb76
taZZodifErq1anx3IyLxnnkb34YE37Xhqj96S9wfN95/eE/0aLXgt7Xmo+CBwdek
K/WqwS6twKCfbNl4DZM6U9r+vKwd5CkdcVmMmRHnt444UvvYAqLNTgZFa/SA3EmY
w0drvkBPlksa/B5RkdHlzwLB4BJi+fM4djX3F7C5rBoqU9wDNBMrV21QDnKqgwgO
JntG7OPAsHATv0Gyn99oGWb7EeiVjnjvnPLLKjQDC7BTQmvMHexELEn9A+q81KVl
89gHSvh/XFKz472Oc//reuFexVc+a9ZTXid0Sm23L7w4xUJw0Wb5MGdCm9vRBSEg
T4CY6qny6mRpx2aDV3syddk9Nwet6tW/tT9vZpk2sGQDDSWxQ4gh//sScsdU8l5M
p6PQIu7dqrGqYEeXRP8rqybLhdbbNRAuMdcHkAWhvF10iGLJzWIJdFxfeNJhiVpQ
GgUqfa3uKVu6akay2Lh0ycJ3MDNCuePUE2Hg3X5pwRjr3LtiBJfwZSb1KhHQY3H7
z+tpXVcZFMNPbJRX1YPDRKkIaoMl3OF5bGgshHdtSLQ0LdnwYYSBfQut2JqIXb09
K06VLzrAXv65IPjFkJitu36hRVdLsDm/cR2K7+m3tHKz++z5he3/fcis+8uO8bGF
u8/KNgVCj1SZYqRroATBExYgB9+qIrBkcJVy6K08bBorH28HRVhcS+EGUwmt8ORN
yYlU/ZjBnRfVTpsB+JH1vR3tlhXDIEqtbSHzyGO8977kxCKQcYMZBif6cIqRkDW5
CwIfknEDQlq1kAD+C1NB3BIzeKe4OI3j4eMv1mlJBpnSr2lkG2ZTda8IPPLhrV21
gqYvjuiQ9RyV3IfpUjafW9Wvy06Tqm46shtM84gPnCU58JtJm2avt+pMRkYqMN94
Z8m4SYDpIwhsDxgo9kO48UMLLOtPdOHr7S6mOHOigrVIDvxGN2i2RjGT/ecYe+yq
jbEbGRRKm/UVBi5efkocxEp8j9BhEmD61rqSH0Uqdqtp1ghZHZzUreaB5H1OByhS
C5l9pbNYWAeKbRd2Qq59F+j1SeJcZt1ymfsoar9nfNWqxUGjj6L5yzsN0BNDcfmz
bkGFJLOMtGyZREl30l1za5Qijc6d973QgiqinGzx2Yus++pgALqTknVTfeMNZU6G
Z6lzlNJS4qBRftEwIAGrGPDhRjD8kRasBZZ8Ve0x+961An0yAlfwflsZorJXojku
ZBePDmVuK8beFkanYMf9jCuXyyBBInUH8zIWYHkfoRyf9gnpWP266Y/+qCB3fJ0H
UvofVWwZ5fNt2DLWdQKiXXBAlnIHEMO9hjmuQLMJbnDlIi/x61dZGiQ5gY7kIb6h
76F7KyteJnn5tPos5h6R8jUveglF/z5naUFLJN6V7wxiVv+6H2nKFPDi1aNA4UNM
g1CySMBcct+778NbMdrx+Pw+CzbaDj5qbhq/MS/XV6YEbYY/H/OfG59IO45rAld0
XRki3/bEhZLRVZCTakG/Ft9kUDbpR/Dxm+vn2Y3mckr40aBaSPURS/DAYkGO9x8p
EUEXGFhxbbfMzBAApuEVsXA1Q5jCasteY/rEwOKeyNVEefbMsClxVsWYykBbbKOB
KlUg9Em03m/Fo5kApys6IYJAkeSz4XktVrLzGlnGnf65tzMfWH5/uaww8ZsF6ffd
cQtFyPPJWfBPkMOhejSGaVg8dcL/omgvWUVhNjVKGw6JEuljtSQfZRLVfPRmjr37
Xc178jJdPN0Vgxyqwrl0jATthjK7cMEJbXfkAHOliin8m4NHYDXG+gKnhcjakqFH
ulEFzj1v2zr6u8T0G0qgXWEhbIj73h3v8OOzQOjmBCSZrbSkum+aUmbj3D3fuY1E
+0FdChJOSdep+welynPEuUdzJbzo6PvWgKxUGV/EWEUScgo6wxWSIOpsRXraoCH2
T/FeJ9CRNMcEjWN4Lo3WocdKMRRQvTIJJ185i8Wj3K6SOGH4vdiY+4ULUsgsEbaB
/b/MI/a9HEvr65CCePbLlxiSWEUI+ngWpca4QHVmdzJgz01WjUtifG4bNLY4zMCP
3699l8PbxeuNUol+T07usQmeiq4dHPKJCeF8+//h1yX6TMG7bqnJO8LOXi8b9hZg
HQVGt75O3mxUDwfUMX9HWK4nKy+pgTHM9i7cOap0Jhh6T9kOH87cb6eqYunW4uPZ
WxpU6JFS1pKghpi52K7+0waSyV/Z5831qifoqtC6YSQl70Jz8V3gAJJ72o2J/TCj
OB/OB2rzcQU2JkMoH2Zjfe8CpaqoKPJZ+VkmFb3QeyLYzWwYsArBtdKgykJfonxu
ltOHT3d7WCLZW9gxBswZr3o9BJ3AJ+T+RXRk3Q+5n9Wi/nHINiiGim+RKmFWi+go
02n0DcAxACguD/SPnmnPMmsbwC8uWXJXu5olmdn2rxIJsB7AatBLU67O/c6Do+i0
krTilNW7JfTfwNUO3pxpg04+q8Vm6JepAjpGqszTgkoQKVa1Du2HoPqRQvrL9NXE
EjtiU2nk6pTSUkZiIl5vGlRfaKnd0tWGRiZ0edTu+GKJ1WTTgkcSUufz96Uchmo+
puxZiM4yxlp6R3BYvJIbZDf7/x3iATZQOZSvmlD5ay2VTHSjvHRJ4qO0OTT1ihB1
CLF2Q8cqsBgYrZlcYBldkvM41R4vTk7ytgArTyuCybzLgKWu77esSHYPjek7NEGJ
LMZH6e0hg7q5rrAFtTHLcuovBdRNKZczaOLShO+njZde2xSAUMnmwZOjUc2LjiRi
fVcJmhsHqFOrTL/wOAkdoptCKWv/HEevcILjFA/VshQeErwfowhMz6QwHveBGRiA
tUhdaLr6yJxiiuwpn0GJ527FSgQ4NCHjPe7hAU9YnJsEqhX6c/f6JPAx+ScONFjC
b4lDiXwXiMrj7P5xUJhA6010hpyj7Zcybz5JWnDNeIToFEr63dpREoq6ZidY+lGh
CK82KmFeMvWLMdIozOapRas/9Ns2FVJJMLixTLpKBbZC2jvXwEtI9WFh5r0B6A9W
gBT6XKHL912PA8ObB8kdziYblWtw3kmPSU+q6MYTKasnZXzg5BF1OPJPCHvdV87K
KKbvKp4oSHNP8IKanhgsLjrMTJL45ta1iCJTOwhxrFLiN+duqN5V+yLzy9o6RnlT
Z3hqNLwYJCADz2sfhI/phL6hkOW//fD2ut117HP8rR1Fax+O06Q5sbi2mQDKdQG+
xdQURE3VoADt17skX9ozGY8fidGYelRYoRWVHURnyIFF4/yVDdXomTNEY4dXdhF0
wRrFFdCDb/ZLRfEsp5HYDwwyNO1YIbqsVDCY+vAEAozQLjB78tTEkoFOI9mIZLCP
/9nOv/HGcC+840973ywZyVC/h2aybnpNYxDvzkG0EODm3EL4/LFIHAYxLjEkrWeN
O1D3pQyoYu5r3I8Tw4RAQcmUNzk8SweF/vVUnvtCP+VXJkF7wuAKxXxQcoXm1y4d
mTY+tZ769BwffHXXlyjOf3/xxSLqQ9aVKDanijJHYyeGchsksdw90CQAPFwiKxgO
UIUDN7d9J63IYpB3w/w7sJkOdsZMdMVFFcwEhFBX4BOv0NUFyJZVNI+DuISYP296
Ibr1mk2rxKz/uue++NSjR5BQqR6u5Ld+HT8tGFEjyfolxijnBI+qsAQlwjQamLDK
1S2DPQAgV56WaKhOv/LHoS8tdc9oz54GiGbX9D218CEHqPPfvJDAizcNkpycAzOt
vMucA1VH+xXR9bmbw61vvIgTibZi9QBFPdBoWevfSP0pkOXCtW5Ap+KM7tvGwTWe
CXipR/aLDVYeeAjt9ntqjJRjVBBHpClsOECeQKqMMxAg+h1fVHjqcdLAoMVRzrv3
OW5cmCKMmmFqXksatEHj9Dt/QMvzdbWkqf3qDFyjyXFGql3t8rl+SPr8K2Ieixo3
0NJFbAcFVwX7DLghEy25vGGQZ5Uw2csGAdxyLhPi6kM8DcCyNzjyn8Ad06m0/s/a
jzLLd4wW1/blVt9myKdqzBAOAtVniswRse3lTrT+b4wrbe3uu9e/MEgGdvnJHnNj
EVrN71ymQShM1uTYaVLT4PtbymrxKYrvEFR0aE5ZvleYMAT6JkGvKMuxWYkWO7Ws
lqEau3mwCRQIsi9Uue1uCs+AOBnW1h5S3gzYXNQcJG1gLP4TYXrLOZvhOU3m9kOm
NYmZMceQ7DDAYjcJcMYugJh8mwPF8IBUiPFeG1Gytd+4kTuoME7mH8Bn1ceEt+oW
KU6IrMOaTXbBlvV5VIMx3Ah5cMSe6UdRtOmDw7VwuvLpGNo0DKER/7S1dP5SK9NB
MqR2/y4Y6xihqjH1r+jDtabV4IEA648j06fm87oESJ2lIqalEAXjBOJV2wKBGNJ7
041JXi2d/DOUNG9dH7VzsNNu19rdNs3VUembLTWE58oG/UP298+BZp2D1eDLaYok
Q8fNEDWcuAKpKxnamQzrIWg3EWvGR/lRYJ6XKJjbKtp0CD5Yq/6ZD7GlHEhMUyzL
hrZFadM1s0BSJfrwQ16PQRQ0mIa1wpUaeCBggmb//+Tgftf1HYOhtq+sxSZfcr50
wCdSwykqZWdNOYmiEkJTuGBWjNAwDBUe+qLXUAy0X9y4VtNwgzlgH1T6BaT5cSvx
tbstLTPYFVmfaR+di6999YR4kZRyMOpOUOZLnOMNemolXWPuo0anLJhcseOzRl3x
o219LCBsqY3a73+ofojeYduffoiIar7+9k9TYUPHASj3hbSAGUrA6Apv9gJWOnQH
P+GA6CRNhecxu0PQtACzhdeLwZ+N+eKzfWYHdAGTKD7ooE00EXHxyFoXI+xPDH2A
J9W2uuC+lwIN1XO//J4rn82wQwf4V+ImZpG6nduIS6WuL5k6A4TpHvCySsyrWB/C
roPdATkkezguX2CkKaGWPCs5W+kpu5Q5AvAokF7l9mfJVWUs6M6XZJ70NNrlFrkH
aEQ83UQtKa+Q0jlaCOE6NwLQmJJkbacMLTnOJcAfOnRndglga7zV9if68Xiq5oL+
FRr7mcv5i6yanojUjS6yZsfpPYP9mKMIKYrLkSNZ6KCiFb2c5d8sUyma9XMiywU+
O9s+XpBYwMRx+S/yEHSJIs3L06npywladqaUIJm5UoaNASWHMcFvhQ+noHSfYtJ+
LLMmGZtPq2DZCqPlseNPiFIJ/0gE4FVQ2kAXxAjY23jU+/OLIISf2g3tXeY5vhcV
JdQrhhEVGmSZjWUI/Uib9YRtc+5Py2q5AzAPTm/TWS05jxb58ZAMgaK9C1qL8ewt
F7jOutfXpsSgkxPZ8IyHzb0BteMUOHVCtSyyH7g6BF+b0hMlhhG41ts3HJsR8mER
HzB0QaVHKX+YfUhG/tZkc5yGV+2w3fvDkIJXqxn6HRs3Jw+R7YSBMcpZyUt5AEU+
mkS170KpO7tB22c88CvCvVJDWdacS/mHkpHbYfmlcaOS0KTEeylzcYwhsl2aWZUv
WGc6zsPEco9LGeNFuuKYSgJBQc+z1Fj2ekKbzTpyeiOabGxyU9X/NN+XT6K+/RIj
79tb/t2fOniB25syOQ57aeq7Xjm3KcB4KIM6U92HU2Pt9lqAwhC5wGNy+Ej0Wgyk
srv2pdmeO1P6Nq0RFSD6kdF1YulSZnTxstzTVMNL9VVRXKiHfopn0Mep550MSdNC
OjSAtYtPrTNets9iS2FC+JH+rqg0LshPYpQhwKQWP7RszIzsEZz5OWci8GA+ALyl
n7fmpbBc9c18nKL9FB4KhUBR+/opS7IGJJXU244Wa60Jz+FulqrTGTny1zk1Op4O
9rxpfCuq7oBZkV/wXcCRJUHpD+H1UegmXWQ3glR24mho4frclG+G4Z8Oad8imCfF
lzYyNzBhfezjLYgs68leFLO/F6KL2W3HyyfRHmSFGQdaHAdVwCCAmqNPFlOhJ7y4
4qnTIuZlGR7r+Y7I2QJBr0IOo2BF6MsvlaOLips/gw9yiJ0lrWyFr5SYrPoCBRgk
fZcWcZmvn7ZFdJfGzuiNc0BanIle1sGkcOPIMPAzTEKsByd8TbFfwYekCJxjwaaS
tcZ6TZtTs6IBFVRGbu4cVx7sh/5V54+7vN7I3WtsGm07MG0TuluaZW3eV58Bn0od
KKORM13dd843B9Vq42XQ/uwCHYg2KT3WXLxlGVElmj8SKjVRYHJ/UxedghzL9Tnh
Ar66pmAqWRcsPZnl7ASyCB4GWRW1DE6/VqhAiICwr7Off3Ey3pRpr7Eu2v49fWny
6JXClyaI/G3flBRv7rE9M/zPCRUfkL9LpuIrlmQNRZyntKgSLvF1yTHU8chl+Rh/
z5Vey64HOz/Tay0THQa9Bfr+kyKZTVvFBwYHRMyYCvA0+TmcsukBGV1g2qQm5X/V
7kGPBT/qnkCvZ53nEKiADu/C5FrB6VvaKQRRwe6060g1jV8zHMvyW9bMtTpTNzox
sz98J6+gDfXB5SnAAhJgEaS3TaHwZ2oKatWvv5ZRiNu2/7Dr1JjN63J/QbvTH3cS
+P1rlHRn9Orbk62OsUrQfo+0mM9JdDvMcQEDldfgiTmbHZX3+yjVTO8qyMUMawDs
f6KJnaSVBlRfFDKjCa0SP/A27m3jBQwYdwZ2S/JZ6+Bjv/b5btvHE3s2CJ5oeeVe
5fuUU2Cj9DM7cBXliytzk1u0O8jiFUZG0y+8eD395SjyNr1FGBDnky/XTteLMU1J
k09N2DLvU1rgLzBpCu61fN91uvgfq3jtPTRQKvsQtDXisEzWmn0qMNyuWJD81Bpe
GQqkC0bQJLSfhtr382isfZ2jMHRv4rIo0OGn47F4dIBx50d/cXAre+E/j8WSeA6+
LNNaKIsjYDOCWtZywUMGL7CEWGKKCyLX/7V8ftdW2obYsIRm8R5SgcDnlaQ+NZHq
2CLFkDKiL+Pqjfn6nNHx/2VUV93VLtIoZWWNnddqJV6EcHP64KzthIOQVc11i84D
vwW+fLBIlT2zHBqpoIxVEqLWYWcwrFxrcPrNJuwJKxl12HPV373OWyk0L83kSNIo
8R9HpciywYSBXdLfpJ9IXsU6yXUctWwQ1mzkhGZ8PnteUkYsClxXXYGDmDWJCbws
Y63VkXCbXMglbIsz1zOYSt2WxDdmEszLr2vaLwF6ZVHNN4kHEFWDJZqpeF6bYAiE
bNZC/AB8EWS/EXS/7qgNxAeOjpeRGert4AtBatUmc9ILFXHXsHmd3sICMrOtR7O8
DvUqNphs5cgMQaTlHOlHPMxd+/UycrEVnx8b+RwgMOsm/DsN2BI8f62j+4FX+eBh
z1XgxH+HhfHkZt8C8BTwBQ==
`pragma protect end_protected
