// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Wed Jun 18 04:07:52 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
VQ2U4vVwGozcerS6CIQ8XI50uL6IPihjdl76FZUmRedIWdeKmthh8IL6iZcC6kMQ
R0u0kngFV5tVBjGxett3b7pJBFGqETJptuxrnWJypIGefcXfhRL67xvaSWI/BtyM
KjfT2tBbcDdbBsex74EQhq5HKrpRjDcs4so0G3I6hog=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9280)
wG8JaDMmc146u9DM8+9gIM4TOfD4wEm9GtI2XDLPZbjLjTVDTz7eNqqlc+4I1AOx
ZyjiXg0CYvkv/tBBKCYoCpcqoah0u7oU4WyteMsUYm1K5ABkZyVJJH5Yc7yLLuEn
C/waS3klu579/yOpuQuD2XNxQgmwC/M3aja4Irgkd+V1/1rn0PWrMpUeDlG5LKnD
HHkaIum1CzcCIAX+9JdTv6aEiprcmY5U0FV4PgnSFLE738H5efm9TPlOQzn0LvBW
Nkbw19jCl3yLQ+bjhKfooiE0f3KFtkY+3EUs+eBPCSSiy7DHbTWA/esk+WggFiQ4
LX29MYlSSz1sd7eClWdl/y0kiYBIYtaHSZqJo4X/TLPiMfsS20F+h115uD15T40D
5K2oFEgtkNx2x/X2Uzdpxh/wSJJri7Z/OM6dtTbPmcc99jmUS1gNlLym4yRvAumJ
z57JORV35ZUhkz+fX3Zt9ATBuNfyYkjy7aR8eXp2EIfRHTNfvNbdHSut6nsSAlpI
09O8RUui3i/iW+iU2r0N7oa5MHVDBZPBZ6ql0EPbVB5v5XaO1w1Is7uwJO9Ww8hB
N0tNH48rNi/D0Xhti8JBtFJQcIITarJBatmbNAzLw2atm553gFz3yFFgDCWfxz5+
w35M6MZRzGkXc9eYXG8Q8DtVExqicaf5JF9pzVoz5e6WgRkBVCsN0VX+INrbzQDw
StfeNPO1vl3KjzK2CmgBm4f22QZSnF9UmGLnUEhXChBPgklZ5Fe62feaxNR3JZxJ
B7xfrVWQz0HhfkK6lqbVGFbh7rvpvHJ5HVDJ4W4S2SaNnmzpcLXNgqAHSIVFU44P
VKcZLyG92ic77/YvvAMwr+Ea0q1MYnmLLZ4vvJdElx453FAvqp79htT/q6tEyIW+
/wQT/JhN0Uf5W2qbqLTlhXw8KfVEEtj0fdxzjXH7YDIYxhs2Qso7X4ckuwL6ci8l
YrAPNejRmLin/iiDeT0eWf0u833tpUSMlCMUkPYNbeJBzMFrCwHFlMgCHA+S8EJo
8rO1YcvRYB0AMIDw9byuJttOWgxrbpw8gGpv108PnVKxGoxT39tB4Q5bOYqdI8rG
tFORrHhzYzI1Oj8oagOBXO4RHn1QdXprizwgkMrbkttGFUg2gVvEpWduaxqnRFoX
ai5PAOIBwPNFmJRtjcJWpnqfxdJ9/2iGwtCoF6GYZvqqnWsSFJ0UnRcPuR5nsNU8
6athYMLQy1WbnAi3MWgekqDDT5yG4IC9VKdUSVIoPNwe125d1+Ci9vt4sjXZ5AZ2
yd2PEMdgPy8+Eh7EXv6t0cibdyIMdPcswatObtIugv41YZmDpKjwuhtrC6U/TcaY
MAvh9v85L/QjFK/mhGOmPctevBktNcowOQ5wh6kXTOzi0CDOUH0gHH3wLQaoP8HD
vxa4QxpkN8bRsXfQaTRDhLf0RJUOz1qaYlUgSVzXeGBpGhZOykxco64yCWGkL77c
50rBgxDpteV5ZIsRulBGXOdq9z7vlghPBz7Fov2eKudppPUqc3AAnkNDtqbn97pq
48OZQbZaZ3UwykYNrsoFtL7lxJ7N9KTsORQmiWsbyQK3uHbSiL/BTPh5f7cnVu6Q
XIThRjeSLDdvdgZzStfTnm1pvHuO+kjq3djZ1H2APpytxFsqraACiKmlebhS87kK
oGZ6Ovk7lvcgnIVtVqtnk4R1kqHMWlzQQdi0M01KcNa50oDETiujirw9I0BMgdEq
/3wHHOQtS87wWN1Fum5JZ190dlxGY3Vnafj37IJmaDDfgPlcK4KBqva8yN3oAdXh
DrM/ta9BlT9gHVx47y/25aBb/GMikzX8NkjmpFCvuUsOUtAAPdFslaUuEXR8bFGh
y+wbL7C3Gc3Trdd//HhxkbWG0NwRn694yPcYp1q5lJskhU+4KqKaZB+E9fyicUUr
2WpkBSADXqaEU7JFEqH6Cx8kx2LlH3lwj8y6BIIM6UJDhGwB8Bb1fdF2llgpGlZG
EVp5Cjy8pxtGATtNualmOtPliUcWNHt0Vw4KZ0X+FI2L3b/uXURHHMzz8MeZWjPb
88OE20EIWYTbJlOFUvdH8mcAFQ23/pcihLt4c6Tep6zwC8zi+PY9n9NNsGPYbbDw
HYf4YMgIFxjccwuROXMCn2QN6x//940JA1FQNvlVHy3AoK61suYjgiYJjerk7xCw
r6FUAYLQeeH/UGhBY0yWOEa84j0RqHzFEGaPu1b4r+0CXekYnGmR2m2k/N+ovI05
8mty1LyPLYju6agkqdMSZ6nc9lzfdDphO46I6rlDDc4h+Lz+XqG5FE+cBxKPpLsC
hntCHluBZngcgduOU0Cd09Lj80MsrRs+vYnr69erEo95CQbITkKo8KWNn1SHgIgQ
T2t/XkVbtCad2StrHb6SW+Xob9xMbbRBgU1aMo+RIbXwj5deFLjdnUHRxNnv/q3+
/0ndwb5hmT+yiTswkhK8eebFqa6UBcLoH/7Vltyi6K3eKc87nOdzc9vuEhYo3R+w
6Lx/FKwbMRdn07r7iQaEEU9nGa/4M6qxM2A9eBlL2FobMGXJCYWnk4sL31FyV3E+
niWVlNtUOCAH/p9xhYE4JXaDzISsQnNDogwsXTssjVe3R3UdXqWfQMjSPuskxwVF
/6GSqbUIagX1eHaQd/JyqW8DX0mCtJijGt9OjHo9uDiSMAs0rCCk8hdEhaaBoCKT
/beRDc5YgJDd2aRSlMniQoTrs7q+Fec2gyJ/0Ct6jgBB2QHu7BoS4rfeEH9OElcF
jfv+beX0j8PqlvSjjE2TjKGLCCeApCp4vbI8rNGfDADXX0CIZMFLV0jK0lt+HpW6
iU6khacIPUexE7emf4mjfYGQSdCb2rhqgEs5vp5+qBQlF/uvarJy3f/uT3DEkKGQ
Ml/1KylIqMvYfMnvU4qlZUdwV1dCYxWK7HJFvp5GWBZMPA9thrmBBq7+vrt7hFUV
Ioht23yTpzoyutrzSFtLWJKxyauNk+OTV8CzHOihAVR1WfWBslWLpSCZ4DD8NED0
Hrtodf+FM4M/6YCloFBJCRQ15OnFqaszXxYOs/V6nKKuunGyTeheeYJfjmxyWVFh
FKLpH+b6wKzR6+RkZ8LdvBjQ3HkEuuZ5ftGBDS8NhJiwtuL0Zo3G8Dd/WcUvtbOW
KSYB8AVm3Z6AzDv9x5zEdL8zwvvt8Xz3PQP9IKOhd/Bnr/78ONmjLYJulzuQo0aN
D0bpcExEsDK7GmnbjImGU6EZY/+vpim7p2eRyBvIgo+Dz80WJa/Jz8a5+Ex1ZM3T
aLVd+XK/8tm3yKRciwZLE7f4Ls3IRu6SS753DtbHU3gj92VmutgkOmpuadbocknd
1TCB+6t4+aCAmc4ENUoM644Dh1/rHlRTpcT1HWNOp6oKsOTRfG0S4bBrSxqzMXmK
P7G6sLW4ZDq3mH48NYq6ldmo9sojZLXBvROmd5F5ubDT2fJpsEquyK4O38oRLqVc
Pcu0ePs591puRIE3ITEz68ouWoP3ZZZMHWkGJWyBtseNdLmqsg88zNIJX8ykEqVS
3fZ600l6SGE5P0eYOFBouwtM2UR45eKNxfIIi1JfrcHC50WXos9mmtRaF1aMCPyi
2vd/XGLjKSqzTNjl3g6gIBm0PYIDjzQzPmZ2c3Y2fly4J5oRNmrb/j96JRIoVtUU
jdpgIp/fWwwmZ1NeEelcPgFFtMFVavF04GxAZGWfBExcH0pEr+jMGOCgn/DYU2kI
XwKyMbH1MGdChfQcgQtGVmPpD7DiVcVDeRXsH0wo+V1jlh0G9VdOMPM0Sf9D4qIO
MRkw7rIhioK3MSM3nMMza+PPQlIhh9Ebt0AScJmrd2cXmhSCBKnyzYRsKV0XAKG0
C4lqUssy6y0uwcFnuZ9YBCTYRar6v4WML52u+LlhWQzfBJPndcRDa/hKjbD2Esq+
wKOPe4KlTS5lFkhEsbUP50P3JTPuGFvOSEzWYTpF2hM4nXyI0z94emKxJg0+fNd1
PVA0SOBoLgsRSZRY0h5+LEGRqrwNOJLsG+tJWwFTUI3fBUHm4adkP2IwJKk29Io9
o7oAz7FajWcNNDLIP73271KhObjDni/4z6dFqZuTpn+54CbhttpELQ4IDxqw2RTn
AGY3aNIU27hrJwfyzhCMHz7SxCsM8wOYg2JbdGWmz5xtuFaj9gHaldwPFedM2Jdz
dtVkNuZDfw6O9OQ1T6B96cKz897sbl75/9n7/BEx+NFrQvgtMVm2Rgez8XzhYy3K
PgCI1uA5Cj3r0w3TrTQLi01TGFw5spTiHupPMZL6XcbuGIFSOOS4tjp+gBe0Cjh4
xdnAb5cwTTpxmVRjVni5iadh1moHXLo3m65FHKvec6f3YJTTpwoHlnVA26Ii9l4u
mdLF1Aa9kL87fIVlnJrBLI/njlN/4yC1aUSXpAk+RBU2gm8b+YVXWQvaSqfA2XBx
5jMxHWk/dsbiYk2RmMB8ZRRwULbz73CwQy8h0bgCJ7hR0mxUcA2yUbR9bsaSG/bj
xinMSx2Tr5sbzHQ489xqW7tIgXCSZNgi6eovcqS40vF9JRT1tbZ4IfDLrVw2l26m
4UFrC+Md8lX1LZ8802+2yuUdBG3sTZiXp6CGpukq9uTqryPtk1VLI3Hvfbxd4RxK
IxbGJfNXmN2wjwPqRpMGKVtKBNIb0hFpLI8BJE/o0ytFJJGXG3eoIn58cjukbF69
jzQm5nOsnArnE/cPkSkAnLpUG2ed9KD6hosy/5U/2n3H1fnQ0m+OF+P4T/DuKm8m
9zwb5wEhbPi9S3Gr97gPOH1Z7GYlIS2HjfLn5pZwpViy9kXBy9qyLqBo0RtNVQ5R
4vhJJXw/zm4xBg3v/SqTuqw6QmIytPDVtEyaxMkQ+K7Sr47IiWoy3W3nOcslLZlw
JJ7+go+5kZl5H5Pge6Vad4hhbpx8VMK3pg9mFHMnJMsCdp09hg/oBAWQP1N3mLvE
kCMXfUd/0yhRW3ChsRuQifJITFoIvHshrsewKmjJKIozrWmIB1wWvaO/TaWFBlPM
v993wMHva2pRVrjIU4cfIxFpH71it2I6qzlwQBE6R2F1wmZCv6SBdgpJ7oMpCSAT
kLV6QVotCRJSJIA2P5stVokvj57+0Eb/zPDoH4KUJvAOak+vphN+XKjW8W1ZOVZQ
4XbgY6YvuJDeTJNsyDkZOt60Qdkr7X7DB7w3Zl6+S8GWmsb0ZfOOWr4L2pJ0gnfG
6ghpZlAsneEQ3G4+jRGgNHIFMWjIY27OepKvOi91sk59ju3RVWE+UVsKY2XfWbHN
kIA3nOgS3pLZMtZHGB71MH3RS9w1ayVMeMIpjb9gA1yks0gpHX/VRCUFDdV/FskB
wxcewXXfqmwhtQKhppZvu0R843rqPHhITM121vrJHChsUC2tKFsY5+Blav8WkEAt
ccfUc0S5K5YiR3TzZx9+xlL6oHDuYYWy4iJ7YalhYUVLw5QGH/FgzuhfryTteGDV
OEPKOYG9jY1iUjuZx2/py+qX21jlkh8jMLLcmrGW9Pe4KClFOTww1CQNsY7DuTPj
w65UtblBbHF6F6iC53srhmKbIniU7QtZExz1fmQXA/e78KPPGH7/WHyqb37dfo9j
+JDeljCTet/QMKddfoXA5VrfBPLMcQ1+PDEZ6vv9ktOwiCDvRXd/KDOAnTHo7+BS
Z2lb9SnXueGs3FWJBH0Um39AD9i3tCUen3Xg2rj3yCJrvOSFlde1lw24MjW/SKrO
NDTzIOG0UdqPnVoIjqdt214SZc4MvL3Ud7Zqt6wffTFa7bmA7brJkOYoIdBqvaxC
kFt83RN/dRJ0GdJtZqzSE9gBw1DOisq5G9x5mBw/wj9feSQOK9t99XmNqYdXl0l0
12Joavp5kt4XgMWQshxVMdst/+pAI4neDawgscrc7WwdxEMSlVZGj6qwDD0AtFh6
RNoksXmEt/ttDiVllR0LkXhN4DArWE7Zmbrn1OQ8wPIQV4i8SZHgllQ/D61AFyBy
LQ8p1iWGMTJyh4rmB3WljFe1KtFPjFdZoXFkrZksRVGNCyZ1KOyqj5P3jKol6Bm/
UugoRVN6J6bXMfMKf21Qzvgsf2CvqUy8zCmjpfUkFvKKiZOSTXfLWLBCtECPEFck
IyykrjKGASptYkGbh3lKf6MkkssiuJqcRf93yA2jKAS4cGCtP5TjCgbc5QRcqZP/
r6YMc1/Y16LYwhfMPbt8o0Dlpxh0IZ5p6EDKKyF/ThFUpkCeYUYQJU/ApzmvPRYz
68qkKkXasx9hiEYeL8FpcGeR4paUAjLr3IJtwRzNuP6TH5MvCe0IMaS/vlG5FeXL
QHBh0eUsjnlOBtiWV92pa9+pcOMJAsslNdn2lxj/2nKCvcDWlPKlYg19Y3GYJsjR
Wt7Pw2b7jPgQwrIdbZEg6lQbdd/OHyJnPaRuaUgORssGdf3G1sED4c6B4WPM310T
T2xTb93iZWncKww7iHPUCyo25h9kQErzQeBjIZruY5Dru/x9ZrKgNB5X0Deu0vvY
gj6hkGw9XEPaN+i8Jt1mzEVdgiYmz77wAiVxa3VSipaNlEcBKVvtDbN+b1x0Arxy
DVhmriOygJvwj1W6hCLhiEO5QvjaLfQ603kObgb244QMEHS2724UEIzajTuRwUYO
MUKOfFBThOcw6hXLT25fFj98k2igwTItgvC6pjtfEfEtGFaqg9KanR93KhQoQblK
TQUafe9o+0+Kqi2A3scZzJwkT3ckV6mNP9F226qOT1fGojRRZBi4SdDqdYH3PqPL
de6jaT/5uIm8Fo1aqSiPFVWBjBA1+SFRpwjRVQSKHx52oT0SmbR9Pd41JPJlgh5L
VgwgU8+bQ4kLrV/ii2OwDYa/trFW5uVLdFl7vw3VUafkqV7JYDnWt8HUlBIZCC/1
elfVmQmNxDoPLCXE2GyYJYPTka9RCKraiSh0GqIGc8CnMmMvyug08Sx9wurYlhol
fnx1K7bnX4Szwiljft1DZAbIoFfdSHUavK/typ1ianucD/8OFwQdVj+ywSJsdR6q
jjNmk8BablZZwus8O7I5v6Vl1pvzM3LGV4cbG8ihxt5m41Lx2CSPc8+9qtKigtxJ
qvvUVZK7JEsXkR+ZcYJvAvPYLaMiBQvHehLWyoVcKJnN/Evrx9mGvfe5LTD4MRlM
yLjNKv9ADqOJWzoDCnljhUhgkpZzGAJYOHstdR9kl8B1GmIj32cb1xpf3tpQwpk7
8r3eW/y6Qf3V8MCV8Jn4Mi2HSNPF1q+85OgQRlO94V2lBKgVMzw9sXcHLDCFdLCV
elsS7SAlS8TKOBcU7pgjgpOpkCt+LDeR8CwMcKQ11g4q4j1anVArEiN2a+LitpQ/
3BepLchG7+1zIqAVoSPK8S1SLOjhdc5xBCUjjUKTqcD4y1LYD446ph7gIdHyXNOw
j/33Mo4xwbZ9IgkZjByIoYyCBCO+ZbMvJ6jD5pEq4y61MwA8Z7wNH3X05gMOGkR2
8Qq/I9/A+xepu8ImKYYaB/X3O6nD833Vcix460FAJl0pqHuvjYiZjBAFQA5iLRne
lxvaVEhtKxrGW5zBrWxrym7Q1cztmhk9bAaTO5ciAMXYsQJmUrBw76nVM7PbXwmK
a2HTONW1Z9svzMaoUij/IWYTmj7t1UiNZ6ysb1PjhuzgNL2ucra8VvYEygf03CXP
GBpH5dA2n+ee8wuKDNCCKyOHLOpMUITm1PpFDtg1xcn7ARmPo/WI7YqZ+UrNjD2M
xuZNvFTxdvKVeMTzzY8dntzJgvDrgC30EakXsitE/YtQPyNV1bdoZYU4bVnNkM3z
HJI5P4JXsv2gjygi9AV8kFrW+ymmhz0WOII0X/m6uaRAuD+zB7qr9FA56FIRSlfB
KP8qMEJMpJGHTXFSOuSuwMH139FIWonwHiWHVrVgOH7HWrLIFv7vsCyARUlVqP1h
+moX0x/Ppl07cz3mnU8HW6iqL/lnrSIj+3JTZ41XQR0PyYT4i4HZ7hGHL5uyyJsk
jFalffK0Hbdq3HWW+D0kGMIqJzAEeCj2j9c88lI5CUIgZERsqxG+i0O7nArW1vdN
tWxJlXlQWuFQwpGsEfM2tMGLrQldFEgrqzS/rLqilDwTtPCfHqKZkMMi5Fty447W
+igPF3E+rDvEy/dj3swQtBIqzSqNSKPY/M4ZnjqCKlug6v9eZna2Ie6eUFO//vw+
bHMFTu60A/zARwZQttk+hIqkOdBVEgxrjzA3maIzTgvi7LI7OLCkyQNDEqEH6RyH
juPIn1iyTP5t5CGKrJU+ZWpA/B9cMtX1DVELJOmDElyxEpbIr96Bolq1VRbMxVpl
NrcGngolDqsgVAHV1Fgsx34WpTD/1qlicvOmPCqLqRCXaSu/gpsoN/4Q+pAx7JnV
VvUY7VdWFzfDjTxIFB9TbliO+HSAGA9bskeotPcR8bkPxMnG6gbyBPOh+LYKF7cN
Gv/jjY0sDC7rgaJM/gAYFr5LaYiJiUI0XXJWxkMar50uz9dGoCkKMPtSLq9MB0Xm
WzZ2Zrs41bQmSPHLqnS9NG/ANeyZ5qjzVYMowoJl7Ez3hOeBa7Sj3kCYoWGikarI
oDwfAUpFU5/vXi/gmnwFoWitVUHrVNY+IbJFo9xOKFFpJFVaD9NnAVzvzE8oIGRS
gHShN7o4vgsKg+k6r4cAuYCf3mH0jDD4XbxMocvUmGy6PlML9F/uva+/krEzjTZt
+0Y1xW2Ff+0LxQ76JbwBSLa6B4tW0FQ4FLpt1ay6aI/52u3NnpQISOXr7BtTCtOd
EVQY/zL9W2ELdUgqGrhKjCxBcCB7cz0aGfA57JzJWJUJfMM9BP/mciHd4BBNe+RE
rF1A/S8qQw1udZUI8hgOb6zShGcX/EWTaD0XcZo6p+C1LrlazDQoWhAX3SxFUfYk
VOdWhTI3u+Je6J0/5op5n61tY2xgl5zapd15BKIi3l1yuqDYKsYb2Yd0CaOdw+2F
fbv12SE1ysm8oatCz2cAfHLVzVa3G+tAS8bgkDaFzoht5QiQAQAFg/wPNDsJBU1D
K5saLu4Ub9a8ahGC2Jb8ph1zmK8TdobApYszkc/pUr8LjxHIP+sakQUVRh743vCO
TTMtbv4/g2f1fRvuOSZve2azZ/mBtZkX+TacnoG7wSvF+8jlLjhfPUekusNjNZ/R
k4RGF77etCa5cnRSoQ4p+byryqjzmQS5KWy7CA32AlF1mShg3uAjHCnOYuoF4A5X
G/jwYbmY+2wAtLKahLSRiJRgV846yVcbzyqyrpFw2PFJENI8a8HyW472xF5VmZXM
19WXm2YkNErHcmiKTb9Q0Nx5Hj9ok1SJu8/oOCRF8IUYwmSx5mAVaLi7Hg6f6gfW
oLEU0Ykj2QYcONeKeFW966rvVyMXUDjlJl5C73AIvPL5rzEfMqxxoFC1pL1zVjD0
519iWpEzZ6s5eLnhRgSUx16jT6Xzzkdlxzy7Z6/kvkRhG9TSTVBbn6XL5ecsk8dB
8GQoXJ8RT/ryODALttMe3TvCIpXvUuamOuets+oPQe9OoB+N80uOPaWGkG37odXJ
NIkR3sXMdSWcDnFHPY4eRmEbRU48q+8o+41FRgfsYdQ6fAvHeiCa0OVyojLDGYO9
ApkAsXrlsDLmzvxSnH+yfmR7nhVPEGsA/juZRocBIV4ypbHelvtz82VaIsgO+SIS
NHKhj0EZlAbn1Gop7bdCD20yRcsWFV7gf0zg+DJhSQhtqJ7laNyQI5nAAjvTRM/q
VwqRLa5KBG6BI6bbYxifWldBqFszRBTCv+DzV0RhGMqljSfuHJ+BHM+FEmFUZt19
moEijv+ed4nCClv7zCxrIRBLPSv/DAPD1fdE54ZZRx28Y3kiAhjVYYYtG0axH/AD
zCpGjVhNYX61IcweUYNKnOKit6rlBwYEMLKQoQfnl14dL3oh/Jvq7BuIhg69yUR3
nZP059H/NLpqNKkC0LJaopEsJ8tLlZqczPhmJIdWEdcV2WABasrG40XesgeWPovU
M9/Ef6bFjvTbvFwyhoLan2x6SVwMC7AOfHuNotVXJ5vvP2QBsTKetpGzLLAlQww5
Kn3mYbxJPczMA+NIPB6u5fEndYukbO7p05XpEaW82XpKwHMelxdcjFAuF3KRxysw
0BBTPOoz/w/1n5dB7uRi5zHG0OQF161iBVmbzFCOAtFU5uzgQTEthXBrEXxK4tuV
HP6NCuXWCVy+tvjeTbYxfS+mWlRJoySWVI354jxHYfl5KafuRPEGpWviOeoqoogn
kzGHqYm5ky+jc60NPMSnLBuaY0UUB6ljnP//xCF1gKZvVCZF+gpxCeShiVIM+exD
wffGAeshxF2GzQ7VzlT/0sYBoULORjUQNduI6qFqIY8wk1vHq1liu24yLWCLDjZe
iMqeZcP3XvQoew9ZhynN5cAirUKnpRx/trhcWSGYTn+jFb7Uvl6FiYPN+j0uNXLy
dmOUXBmS3Hylw49wrlO+4GHdvujFfziKR/WYlcpceAtvfdbFSv3nkc4Eqw3jVcdb
hnpKhKxvME8BLLibUzgG1VzY5RGelUmLrvWocIvxLdqINGLHPDpMm3FrdDFHSApg
E/gSbmPN4NM03gP1UE1szL+XxcEQJSVtrZuWCmHnmv7Rf159+SUlDhADiqqONUIm
WVL80DA4rbKKNoOV5b4fHSP0xxTQYbtDfuNFVKSYSgCnaWlCc4z+XOXSTiDRISYH
Cqhx0aoHDxfrdHlhojTNNddbkPCkcWcOYDpmM2mT907sgyZv3gAAmG9bHBno0Qo7
ZSJxZaL0OAxFLb0VV4vo4Q6on6+fNRDQg13dhep1F9YkH/8a3feAL4rx8gUBF2Tw
CUKoFeAGlS4HujScbpOWJeGYetVC5ZMzW9MddW57XmNKwnZ9+kZU8s6e4bFwj37e
ru3KeOmJ1V1jBvLGWMukuCSfeZOCk08Wk9aNOjF4wd3N6GQAghYff2TgJg+A1Koa
BUhqPXZpaQYFQTKyIFAvzIOWpvpbL7iLoeEx6muy84n68hLTXUkybBadqhS9LYaH
BTHzYPN6qHswtlzqOuNHlodvUBFWejRlHc5KsBGPZMcAq1y5W3TDDdxGXP+wpucQ
KufB/EEsSKeF4b9RonPn+65RbNpNirGkhpNLuP1iZ5G7NU0Rh0UxoFHLOaoYhuZK
GnCf0Qwa5Vh8hiQL3qU8rhngHiHOSxZUs4pDs8D3twoFD4OIpgioZBdkQZSjekBh
84z9L4CRaU5bdIUxfowZG7GvUbkqyqOo0OANKtqM0lpf76f2zJa03o3atM0vSpW0
KRk6ioOwtUT73iiPN1W+xRijeKh+p0FkzeVwV3IfV+qB+VF58c3atH2a/Flhah/Q
J9oWoqhccvMzg1AiA0UoOw+smmI57sQXxv17p31GrC2yGLrZ8jk2ZNnp00+QuktV
w0M4OehuGanBE3WEXexQYiTt3Yt+O5PgkoOF0/2vHjC1gMISXDbVU9rp/XyBWi5a
UkWIQcTrC+NpJd5lcRJz4EC7Teef3v4MJ5lKWBuCcnLt1PevOVPQ+Ceq7UOIH1nd
OjzMDmXH4XYd0K2JGLz0n36v0Y+LPJU0v0vGDSAGWCspU6J0om4p4vLdLpbRKeuH
ex6xVnrQYNlZ4Hg4b7uvUyeR2AGLHjYgjTFAJuxPEC/N1QA/Dwu9yH38JBa/I2lg
sDsZv0a5h0/ntuWdC+QD3ffJofxCkn5WXk5uQ5Cx7y7S0ZNn/LUhOczSd7ECdyW9
CD9hDV1v03+0IxxaNKpGiStjjKUZID9+62wNlc11NDzB6BD2lZ3SvK1Kidu1h+5d
vxj602vpOCultjRn+vwydV/R11CX9MHbA+1x8KH/nPW4S+myvxLjwSVIJNGqAHik
j4ksR7ZWqh12OC4RTBpEhmHomSU+VCG2ZKf+CtG3POsqioGRrPSh0q8TRNsIaT3e
i9ZuPCnyyUNkhX+qS2EWE31ZXhz37VXC+WFMa/6d5Q6DPi4hw21mOMeyQSJLk0+p
r/4c9aAm9usxYy8yiopmwWNBoNspiFyJfccDC7/SnMUEhe/+UHjO6O58DvIwIrFk
PNMp6okwuvq9kyjp5LOIKeTja+TfOrvuCDSjUvjenLNONz3MAwXbcV24Xc6ugtkp
G76buTXj4TPIDq/GLzEa/lD1ZEJu7b1dYll2L06omsnh4Ks/3BkGsTy0RlIc9gDq
UfldN2lkzCKZ+MzZZ4+ran+JMn8cH5hycQlmhx4MbzHICCIxkVhHD8SBKj/MmL7h
5vWbiNZjvkx0n27pDtQJ4wbtzv+sXvUAV9kpSm5YaleOpPU0LtZ/j8KHNajaI3Qt
tH928TxjJzyijvNtjDQR3UGIAvHF1OzljybeUlLJF75l5qMvG62UcBajLT0EmOFV
7ptOPpiiq6ghOuZE2nCg5ygpNkFVhbWAk7UPEUht/66QigDLtwEyVNxIY2I6vmJu
eYggpBMArpeqp4Sz5qrNSQ==
`pragma protect end_protected
