// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
mUZxeUv5Kud9lI5mOZmhOD+WdcJe25Gzxyandzr70tjcvmVqPlFMUauQUwhHwplD00sD6w8OcETB
RjcSfq+qH46DYRGAiGVqeql4cN/clP5q+vRrOsTRahHx3UdNi1BLT1bs5t3ya38cRosBh4BtgbCm
JHyI1ocGOfG2B6Pnca6I1mFAT9QVTypTwyPLIhZLgrWPR0Z1IL7MMi2SXgurg+n9TfgZREuL6Pbi
wQ47EwwJROky3Ke7w+nRW8o/EAFHB1Z8XkJSfc61T6RcCiG9nQ+Gu0IEm9nY6v2KA4FaKhkrXbrv
lpKwQ84gquSUc5ijHwYHVfO63ob69VCTH40w/g==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
0R+DUBnTcaENpwslzxInMBZL16Co3/KtGR5/S8UpEu3FXMTJgndRBT4sSthssx4xO89qIvu4nK+Y
5dKQyunz2wPzIUOlsERrGJ0d0AVu3y9J79vXzMpU1t6qEJPLO9jXZ4iRz6bFyIPR8LzMB8mePZct
wQ70dDheaMCZpU0SZnk0iR8OWy3ZoWtlsjaE+/GWDH4swnK5d6LM89st4Nx1bh2+V+I6TeP7ydtu
4ZT5CVBwK9odFmFjlOctPAcGaRLf0xb8xVUrf5mwncDGujfVrURSLo43bTW54fZIfqxY41sQLi95
7c37AQWO285XgnuvaoFcQsmPbaNrhsqFjiVP24rpLWzQT580vtpAfB2cX6Q7Dj7m3PjM1W0fIYnI
45IgZfrUcNf75mCKrIj223Mnq0HsECwhp5Ot7/lsccwAIZ/EKHPLDMoX/5j3AN9DKc//lY4GehPS
P8YSj+EwzQD1nbXOs9FLiKCPiVcMnLSdsPepp7bA4z4apc4iAiXrnckROPAWxt8cvAH2ehNiEQsD
qC7KfoffPYnZKmDPQrEkbJY9yzHIm62V/LMIqdS9nstv/Ki6RmF4GGAFaKS8tl59zqIB59GMd361
sEXfQhvCKOe5bQLdvw6RFYs0H9ME5S7E2iBFefsdsg0LI9LWYu388Y5sFh1vRSiIlCOmxWck5C8X
IR0WTnXqgXk2oOVKOo/xHZHBSyw/0Lu7n/WR9BWlSjl6r8AQoV6+gH0EClRGBI1Pml1e5ym9HMO7
Z0G7sd7kDpkJjruEqTv+ovYquW4xJPqp53D23PAWEbXiXS8DLDAlrWFqjR1zYX8iu36cCJL/fQYn
ZEjjlDgobGIU4td2ryHJfTAYQZTVmQ6yC0SQ2SvuwfLXv2Zmy0KRJhgZojmfXO57MDl+In4kfuwx
Inzl6dmLUwbr+Ckcz/0ycTyGRlxhvArgKfMy1b9pcGOTR/x8rTyD+ArXSR/WgUo/KRYaWgv4jKF1
pvOjFCCSJSPKNZC2cgYDD8Mt/rLBuufPvq7knToQcl3Lb6+MdQDL3JDDNVVAIDFpw7Em1RnKLGM8
cyHE+M6UkUNHIu36GgW0b1CU/Af9XgHSOo9I0Wo/qbPGgu5AcxAyWOSSukFPWay9eRymi34+31S+
Jkb2MaWOZYbDKKSlLdgAzsuLiJqkRkaVqM7/gyPOCLvyxu6oMWjSnAXM4u0h+sxkPbXI6O9Tnkht
x/lOvwQhOZBtYQjMRs8i3Ry6lEVMWwKTebv9nnzfxrMYkhMdz8myi2VVCReOXz/8/VZwFkB++W3k
URoI7pN00v40NXmHg2FKT3N5TCg7RGo8LqbGGJYJN2KlAtg2BM0YIjbzmc0AgM1nrWMx0BD83zH5
UucANJ1i/Wrm4FUFe5teGmFUVcE+K7RDVZz+GpFw9aWYkxdQAbCxbhZ/3CubMgTnwuoIASasfwpS
I8agLMhJa0c33IK4mxTaxpPk8LMFV+GWktNuDKqExjhPqfxjQoGKGRApjgt2rd6Uqq+ZTCO+FCWm
AT7O1M2nLywVbJuZFEtXT2awwAUN0R5tiAdHIIBcP7C+ywFPBN3gC/hNx9UuG+JV06g2OmPYLjs6
FUTt3p+IRKwvQovlvCtRdEjHyp+KNETUwrWS+jPohzeYN+Ft6M6hgrtSN/tc6U2w7reV0ZH9jvy9
M2IFb+mxfl+OBVIjOsu9Zuur7lRUOlWDba49o4zmsjkYGibFVmSpRQyBFwxiWdmzyNUI1p01biCa
F7AqixB/MMYpl2DBEM5/PhsX0/KipFgfTY9GhXdDeS9mpy4hLe2Xo+SD4Jk/ZbBMDlcqIPt21JXg
nWystWm45asllNqo2V+8rC8fUMBYRQKmpwsArILQqKrfNGQ4HY8XZcZTGiJxErKsxXTSgJmmRYqT
sJVhvSFsirCClFQT0FURTRsLMJQ3u3oJ6E80FltoRQE31xWDSYTrP5AXoCfLXzhQWmKkhiE+TR/+
64l/FPDwReM45R7i/VcQqFbe4DB3TraTKw4f+iE6JMx9JZ2Yaf/hfOeQ+vbhfBOuN4rNxZKod8ib
dHn/VHT9fBgzpNfT5LATSCTF8Ih55+Tgnw7o5j2PRoXfleFsOFJb7mjb03M/n7SHRZl0toRgXGcJ
0xqHWCnc+yW+EEDQFVEolr4FoGM0jywggfcpMjOW5KAEDlwInew/CuHx4JHmigYI9Jh3T97lc0KQ
VkAMlSH5GNhyukW3md1Hq6CEkAy4K5DkoTswlLAxbFfc3xhFNKoOjchoefjbyWn16+LmXGFxO+dx
59piWyr3xqIEWjVop6wPro80KmNC9fZPZINhUm8nDc0UddSouL2HBh3a8qlsInRQX6GuT70xDM0V
1CBrqCEsNyCnVVHCjN4KjgSgEwQMXSmKDQd7npaqjlEsWzeDyzCti7Zs4/dgk8rOUszxHzbYOWRV
kC2aVrXDP4NuwsfvYJkfN0tCM37mqZmT2Fd12UI8taqosbfWexPx/cCFNPB4dR7ZCY8Zr8x8FNO8
V4HKR5jyy8IbvZLf9rD7Je0J7bZfME3RnwfQpExpUko3VYWFjxIDgjl9raS6sQxAAk+5cu9vkvPF
Rkbu93/iXmY6FTMxyYiiROCuau7FpKTMdO7ew2AOhHK+i2LvVG1Jj805aTW1rRjT1m3xLupvvQ+X
VQXmA+l5j9d6F+Fh7+MWVEv65IRR8Kwz2fZrAqb22X7fdJQD0fhjxydqTay/XWJnaNEDCMfvhl4V
YZepRP2nxtSXHyDvOPfOZvOWJYrEeYvu5rmXdNqx+87BdoBpr9+hLqqCCPRPbvHtJR/e0c2ruLbD
nI7OzuA32SJn2zSTapYCklDFuaA1QumKVj4WOWA7pGcSeq4hllUCsy9SfWlkTWOBuiCsP6gRx6+z
KUk9bhBBQb4JHFFsVD6fUMOjHGGJn4ME7akHHJZkkdpDBPmDf0sPSmBkKozv3taEvda/WB8RfOPb
AwjgO26vy2cxq6MY+hF+WBZADNtPnZfnaX/mcPcEr6fhto6l3m4rokQrjYW0crbEUAWIUipRaIcA
4jt1bnwmfXTIGu6/toz3SmO1ZpJUghPS/7/GWP6Ub7kLtNy7lT/9ycC3WP379zYBMg/tXKKp+LQt
HBohRqFFLgzd9mMnFmCUScZNZgos8xjZ++OH8li1oXY0JhCvjoKr282RrKvql1UoL2WRmtlSY6Vb
PwzbUU1q4YFonw+2D0kqi41F4xo5wSWORl6r2Ihzc4m/2yKp7j7ADt6w34L8tDVBZ3wfP+ItsPZi
k1PRzZvLqV0hLng0WGe1+t8GE3yB93GDmmM1h2D7cJLqTbdqXj1Hv02/i/VtVfUJALb7vQ8iYWrK
R6iMhUD+6Hz7Rf9oMJqR+rNa6QBJE8JCqWQiIDUnpvYBBfMz94QYn1IstH+gfPgQ4h9IeCn/+7fA
pRvaCaaoghXivtxRZWn6gJ8yHIQi78VRjFxQXRpjPcETfjKF4dyZXfiuhpKMvD/E6hrQHwX6OtU9
YT7tW/z4/bAwx1lU6LpKrUJ771cAArm72ifAK8UixKnU96exHN549ExfCiEF1qrlTplldkq97qv6
LMuc4oeAbEfpiMahG1DSzlYzTfSd2KCKpljGEruwSOoJK7ivrlpoJXXiJjNHJJRbvU2+CeiwCPwY
TR9ync4klQL0S39OdUIzHfr4uVfpf/7I+b5gCvoyiKvfCXbgL4p8KuPQdG7L5+ZTsV3yYAshvenf
IXtll1Ud7Qn7WH3xXtFWYSKDWcjY+teocRMN+DUuJGfxXBZkBIHMPBfEv6dXC5mBcXwTDZ1SzLu2
nJxILk8kYoRxHrTErgyXKV5lJZon3URE+fEpEr2fFfjlQGrGuyLZ7XZFic6fGjFRkheJ9L3EGLXF
F68te/w3JaWxRaN6iUjYisuwMoxrxT7vKZJV8WWrP+anE6L1RIUNnnaS2sD4RriQWKiGfwi8OmRj
iiaCJ/u7Ee5mQp2my5ipxuZ2iTUlj1ejoQiFvU7+lloRhhX+9nAgjy8gCNDdDS4p0d8nawGAeeLj
n6NqgP8BS/O02UwEfu7cf/RNxhvvlrBfPz6RMAeELVi/3Uw+HYwBsjbhXM46/mkIK4IR+cCh0lzC
PrYAcgoPNNcwNbRRj7vebicooeyySWNHkOJAeUgyXVDCifyrp+/nHiYdM3B2JmB+SQNcruGW/4Kd
/4fp8aIuN0kynU/6iiGj2oznUt4CoUySbrCd9fY0FTmj/auw7q3GBtMeXudqAiqyTXEgj4p4vrpn
mSWBSPmU/5f3wDoF7xamPklAsS0xLT1NHi+b/RaD2516AIXsXnzuqQxT0Z1a8V0zZ84+9OWujdq0
6VMloG/cH2Y/TvYhidscGjfSpwzS8IvmSi5JwitKcfeCYLChIStqslR8neimiUJ0mMXyiAnlJnh2
BJtXxvQOG7d2lCs+cgEG4LckuCi9KsdtD2gJnqp1ycuVlwTd5CWKeDXDwZbK1fcYNUCaVR1SfMyU
+UsymxJs+QhqCo2NXGGmAdr7pq99s9n8mNUu7AHbMe1pUulibQUojh3sPY5mGWjdLYZrHGWKJdga
0mBrlfMbBpBaWgZsfAkJSq9tBj/xtd7MYB3Jhnuoaa1E3DfkrArBDZ0SfQKths/f2Em/s1rK75GR
jugLc5agGgtdcdY6EP7GioUQ/O1fAfVcN1Cf6hUATQuBHD46zjG6D5v9yTFiNBFb8s9bW3qonoMI
Q0ufoubAIUcbsqEubPv3GIYdb6mtnCMevWhpMCV1rtHh9eCm+eHjwviPJSl4wDio9j3+A/q0Yj/9
AYINd1jpcBd1J100oJ7MBOdrF+UAeU9T7indQZElrXHwq/uiQkldQzGSAGI4fC/mvDZuU+i2O5Yj
YklTlYsGS2PlrtYmDRLBH/qOwN1ukMg24oaHI94igqovLuH3N7xo4dVGEHxjw1lNQJ+NMgEy4eZk
jzieV8f5rQ1stKCfIuTBic+Zabo1djkjrlG11gmRjV2JJVJlGBUvExx9orlmSCAGFJAzvvtdI49y
5gsH40ddrQIiMI9pPAmsnz77EBETEnwLxqgF8C4MK5EHdzm2SCdb0/Nj6lyZSZpNSnTJ5V9ok5nL
MqWakyfwp7AdYVGF8+WmqiqXNOdg7j57tIQEGovPhnJZgKK1SV/uLra2pdNqHUAEOd0Fcb3VVG5a
oQf+gmvu+BnCH9FJW37oMhPMIXjCAH4cIuFCOYO149P2ZfGQVTqb0og0tIevxWb5Qd2GArPRxdV9
6OjDUCIht42oCnpOOENgQMattmmHHQ+JSArCy7mFLXQDl9DJVphZ8OqdGPIdWCrRqECyGFFx82kO
n+EyLYNhyWZ1up+5OJAV5zAbgx9aQiJr+Z39j6XshcwYvvvLoOD7F4gVVSgmPufYy1NnlsYAEZeK
sQuabT11dx+BV6EFnLLoH14zmiTSp9n0bGLaZvBPiN7nr7B5TJxoSf42DhJx6cx9i+BhcrgmzGPu
EmUI9nXGMM1I1A380czurL/QhCBXxWfoqpKOtQUVH5xfIAUeBLyIzbhI/w1faAh9AdsONjZHhj17
6nrsX4Mk2B4J6FeyWFNkLVpDuodaZbxyU4BcV1EJMBqk5squONSi3Z+arXqpvSs7lh3wm4Nas73r
YKae1ENDxbzb6cOhKmdno9/9fG7K8sEsXhvKbj5L8EaA7pHW3TCu+FsoKA1dD8Ys6uoaZL6YAaTX
jPrsFFg3Sqr2JaQNI4b/AhacsCv5/4x18GaFlfwxKAlzsv0m8vby1EpfXVfL9DewA5auGlDNgxmu
j2M5R7Kr0hCKaGeAjTdIPhuke1nofn7odpqNZZhDuUsdvbFSc0X0TA08Zrx5TtT8qHg4iXcXwni0
AS7K4DxSzrupiT0QJ8eyc1ahLNGkBc6TSdjiceUuYrcgpmhl0tJ7f2YRcDGoNjcu6PZY2sfpRRsH
wvsJ3ma8HjNjnoiSdYMA6k1yAiztn5JLswVp3VpirUTWNqP480HZMsN1OcEaGyF9UolyngBOZiKg
k0MWQodr2pOAZWIa68Gllw4uvxtVSFWTnvp3M6mjd0JmLuDUGxZLEVWaso2uFJKuv/sJp0A/huLn
3dPLAjXGfpVOxVXIDBfe2qnweeqw0ceA5EKOvkgCKE48l+khpQRJpnQ3HpcUeiFfTmtEVEKk0vT1
AQwb5OUl3BS8QUW7lQThTlJ/MjssaUbT0sHw2Yp3CCdAbnRmvHi9rRh7DtgCajWEG+pa/qLLOjqV
bEbmc+dzBsmasNNUIrlN1UBqdwDJc2UPOxcyhwbEwVZEz0srHr7fni/f6UrZAKJRBpivZ+B/UAfp
025im3B1mn+qeif8g79daqQBXkjPwdH7Dz219vPP779i0GV3mFbynER8GTnnpIagxYI63t//ZdG5
SYOmdyIIDEXQ00mZ0wuEi1NHrod0fst1ns+Q/SX8DUSZaQUinprZUgYf2swqc8St3g4WjJ4Nq1MS
uzu1+/Y4Ogc4HEYVIbxr4SRw/MoWB8lqd1oJKE/yJSOu2ZUUBXvzC0cO7gBQ4BNn4FpHuKKp9ihc
ZbabHDjJJnV2e5ATDTKPIAcXPv+9W3ERNTQl2xQ/hDcdhVMNRG9rX+/4vE0PSEl5z+w0OciJbLYW
TT/kcUQEWr65+Oy4J1a63UILIaQhR7ji7qW+EeAB0tAfAbCdPYVgve80J3Pc+ay+pWeo5DODF3m0
KumLHmm8vSBhmndZxYgTnLzuGcP1os9GU7sh7NDdjYfX6SWqZvzxr8lxMXhMMXIQ7PQH2Lwj9Ois
mwtXi0S4Xa/+sNLKEeht86DcygsgQAwxmtw+76tewaMag0mzYI/vrC9VLUDQHgWBoXsxZFyOpSUZ
3GLEPOnek0u9MkkIy0S94Skv1ntzeQvM6phFIHN8jybF90YW/4R9Cx0tE12B/nxfwixmxVhydycn
DYeOWjr42VronvfnsJ8Xnondz8RTWW9GTwGNQau9BZ4aEszHFrKj+SHyUol5+UtHPsBVT5iUrSOc
rcKYw8HYb5kxQqFyKXK31mNpLJZSEgrfhXrSvCFTiMsSx/5maBCoZtM+kQG5yEnXxm7ZVu2T6npV
7kILeQl6CknjTHkkD/MwtfldvLCmvuQT98cR/FTyqg6yWDPf2hky9PgP/6ilJkEFoTYOu33V4QMI
F7b3rIxn8ER1iBj5TT7uCe6MD2fBGmWh3YF7K1IheypClelMtgz0FbzdloUrPeWmRPuTpQYfYVv+
I2HpdoFsCLEa3+OgU7R10XvcrzzI38M/8Jk3LqGv1Z/VGKbOscj57/m5hFJ0QI9rzRV0tzfBV2FK
mtUk4E/hFgFtSXQ1unT4hN4cgtqj92n3CogDUCLTz1qqZsAR0Zl/VXtQ8VvkReqH8pfA5khQhY7u
5JrGd0BTn1k9EZJV7bCTM0tbZvxtg4f3GDJT338xaIa/jXnzZIh3ZaoZj42vTHj//52gUjdGvOhB
9apL31/ro+wE2Qfl4kHevYGbYLpt8S28cyovoSRVqgaDKjvEpttpT43yfuQXQsr6FG3gUp2RxcRe
hzMzz9YvaE3qB5eHtW/YdwegHMXMgCI+/K9gQJ+luLHo5OGuLBJhAaq3FB9YVVYW0KyjSsIRrccz
2Y+evCfuYqjuZgKbn4PjaxoQvO78sVxBxREOOfmvnFlyrOtRNOwGT/8UN5AAdUcjV5BxSTzPCaQ6
7BnyXy23P6QwKtb4C+NPzPoDGMsb51Tv/01e53A8l/lFZmNOlLt/BcA/1/bXkUIbyQvFohdz5801
FAQZGjIbYtyaqb8/W4Lu//RoyUIZb2GmSl/logCSvhTIQqhWNLzR81dHHsrIlMZ+IR92CFtpeZJY
BaC21cgvdPANpLI/T2vdaKkY75hx+VjNvmX+93aJANvw4YX1/cB8RpYUfJFJ62V4H1yiFz+aSVut
06kKs/+MKfyFNdtXvr0AJrd7IcqiB2fsvj17OcZJv+n4Hwqb7/8jdKsTy0JNv1KW3neexf4+UXEm
cQTqxqPJDFFOK3QS0Am3KjQLqDzpfSZTquXiX1WRwx/U/bihpvohgiYZMKF0tvIIcby6XEkHQ5DZ
3j4r2wFMzjek2nTKMKFo+0tqRBvhGFIDFsSLyZzxcn4wdOz2XhtA5g/Cj/qDp82KHqj72BysNTdV
pFWyyWX5wYMBpagHAmbb5d7re+Xkh+YgGUKOu9uiYP4Q1rudxi10ye+6cI0KHII278rG+7UCEVLR
i+7WTR9AM6nciPP8nTbRfNNjbVPy/KmUMd4rWLH+vKJAHKZknvo/JIC0qvt5K3NisEkf43pmxlm/
70GUEhCulj21ejoifU+8IEneeuwbOlXx3kT8ARYNWefnziAL8qGIX+nKdzayws4hC4VzZrVhxslP
hJnVfDfuRuWTty6I0rzvmlF/MOLNyRp72MPiBGYiCLEZtuBFEn1yAOYcWRCBWADDsfHs7AuSL4Zx
o/HFWGA9oQxyjXC0RktUt4bNh3uJR24gM6eTKwHIIdVr3i8A+jGzsTa2Z6nTNcVw2hrZYK4n3OUs
ym+6gccvVp+kmld755rgPI09OqLuIzExf0DuD/5RalkZlBdG90NTW9JZbb0EkeKp6m67Y9AOXEHE
CQfuDvAQAHVr0Aa5S4leG3sxg2huPZqNmjpYeoS/px8gwqBat7l1BOo0fIZH8ZbDxi36jtoQLOT1
ZI4IP6h+PoJr5Lmd+i0M7uRxVK6fJSalOKOAL4S9+8eRg9lipuufIB1eeRdSDTx/sXYmJkDNBkny
s/pnA3sb6kD/TChB2++3+GlCIJvWJGmlMkldvhpvru2sB65he12ALdK7/jMivacJ8jkUsBvKmHBg
zxb53BwW4vrP3J2qjBGeZNg0AMiQUU84x2KHBISNlV96jJa3xT8FjTbpNIyj9KZiDXUP7y6ZCYB/
racit9A2uVrGj6P6V5jpPJriXxr2aJLyI0cuAC7sTalyVOtj9Uw9mC8gtkZqYv7kRzVq+CLI6a8y
RtLHa5wAtSUuK0PU7fB4GCBMoRtG25fNQa6NL/mEvp/W16BbB5PWRpAICmmPyyY23myTdS2VWqAg
nAh4441UgqCLcIwtfmpjjsB+54Zc4TM9Dir3CHrObZF6df2ZTQBdeKS3YKx+v8hCq2uc8eXPm/5s
9grotO1aHNVabpQ23/UyyQnY4sa1+73ygYLyezsOdALpLifoi5sXRKTtqdyFqrHyR8dagKXaG9tC
xBVrlJbn3oeiUhg4oRQUhRVCS5qaXbS86QpnT7LVN1tTvmbOL4gMtqnLydTCq5LanYe609NMkVlh
lF3DbuOjYcKdzhQniOTfXHOWyNBcx/A7iC9qzV/Ufj8KMaetHbS5nPjbQWv3DlU6Cp5hH5yJWSU/
T07cQdqWRg5nuMru9N5TzEjQzZWXzx/pdmAb7bSYHblO8HTDTecJujMGGtv7Wb/V5eV97WeFtGN3
yOaDjiBzpzpm+qLQkj2BW8FgCunSmvBRvGAcAf5zDavr/it6o7lL+OIrzi+zrjiLzPcMKHgg3lZi
2cdLzkZ559GRoUxPCDy9KMcBJmqjSC99710xqz37arhUSu1Z8RXVhNu30Dgs8rHgq3i3Gpmw2knt
LRcxBpyfnOykatJYuet8Dok3Qr/fGbwxkXvcH0G5EXlJtZZiGQQycw2qgOdm98YILcz7w6ygbq3E
DPLcTfKbcNXrDhuvdmLS8S648zLGl0co9Pzu29QjOWgfSdwipXpWYAqAT/HOVvzR2PQzACQm61aP
15FnokPsV4imjE5aRfa8MxIhwtX7rWaiM1GUmo/2k+2HBiVjy/wtgpk9ZvTbEbGuYqZHeVrTe800
XpO5CVn28pN/eFTFFm8tvLiGlTF761SUnVfqPxY4nKuBCvYJUkLyCazS8ZMkf1CLtO9gWeeSHJiR
hd5LyLRLpQuyI6EzJvq4RsFG2MLYQkbb7APFArdt4ytY5SI6iSVVeiD7ELI/LokARPa43Mv4JZFV
w52fsiG8FZznUglMahJAFx3mA0x2gcF5sZvLm3KqOATcDISj2CMy1ujNJe8DReNdh99z+wFTPOUc
90rIMWuekkTAIV7jSsntZZY6qYmJk1hsxMlvnuGiIYObtKrT8QchB9t2llqVmBdfi1g8YRJ2nwdG
4aRz0Xw1Qe/yfY1XP+IQczC8CbPXWIjA/iZtUfIUeRRLQFBLxvQGIhw0+tPgbulvNo65k/HfAZfS
FTU6p9Xp7hyl5b7xXuAgcrsCK4TzT6WSPTKX4p3hUsryx4NCTzToAiK1Gjk2hEfYL5yagdAkS65s
kLLJWz53q4om9483noissQLP4vWijUXIHVM4gTrXSkTj90Y3vVY8675BJuNEsZPSplMwW+A/w1kC
SC1M2Dx75qqVXTc+PTWg9GxdvDFvi/883DUZh15RgaVHbgrGkPIj5ZIHvpecuPef68cd43mgTDxS
Bujzir+O6NHymWytegBoZEe1+WijtpIMdLjntV5h4csEpsRFklBW8VwU9aZDITzxV4ifvOlc2PBD
phtzncCriihxxkvgUti8XFbDK82+x39DN60aNsFAf609rqefh4Nq4l4NCYhaL03rgSJHz6FS3fCq
c1D4/HQ81pXYfW02l7zoopXS//H+dFXB3zrhPvM39swzMHh7KzBt1Nt5fN60prxEoDfCzksrzwlW
6VB9edK9OAtTU/bbOUEAyY8D1rvlwx42/tydbuBwM6Qke8a6kggg8RsojptLSYwA99ySUreOUrrE
IR99+Uw79bSMHuI5eDsYg5wF0lvY4LmuaVT58nMob86OJO8t/IxkL/lGWpI65lBwIJUbLHPme2up
TLX0TRQrm/ERQgRp8O0+ZavxUT9dDOInZq3w35ochE4Fy45U8gHJsPqRwAl20WUatUbBLSwPBBEo
Idh4XapV8oQPfm0K5uhqtATrhzMleurx+Dm7zGIX4PI8zYAGhG0Wkx1OuAYOqmSb/lufJXcJEhiV
CFPEr5jvq8IKMlHyVUqM+rPaTSNKpwpITWNZ420k13A12a35wM8uXXD4roSdBRUBL7cBU2MVP7Fo
8SXJjpOq6L8yoQ5u/Vbqhnr8nknspvvKu6JWBgeomDq6vY/awlHalazoufwzotAIcCvcPMK8BAOw
plrsixLAeIg+IO6vHh9D/xo8Cc87ppmragr8PEvi2yYw840VeblPCjh1I2zSIRHYZjfbVwnxC9xH
ygtuvcnWf49RuFXMUl+WWwyzUOty0nuRVoYMQTP1g1U3LO5pBbdfLBba5MkRveroD/bO6DraIJwe
mqIeS8GNFwXl+hvreIZeNDxDTdFoi1i93Vn7c73vj/Gl4rSWpHcza0UAXWOIrgTAynqbx9o8FX77
JrSgvG1tBMBucJ/UdIUslEXaKRZSBqcgqWmSOeDvNDeZBGiu7U5z0aoiji+Qu4gRAY7vNqMdwKyo
EDpAJW6ic9rGgwpeVFbk9Ky/E+48E+jLntFfz8SXnjCTuxTbkRtb67PSgyCJPwkKp4AtjHTebq0m
KaAUKNfJnfw22IjDWBzvfYeCmZPOeSAQyx5lutZb1XGVG5Ry9+XQS5GOxq+QqZXsZTVA1oMwutKS
tVET76/eiboyLdTNeS2MzK1phxzTLbGmBe/ktK4LF//VvllgvDeXxJGCl0eGzssFnC2zP0U4NKKg
3eBtbp+CtVizzhWcBSkpOF/dL7yp00Umm9i7f59CROU46Y3XU6W8DcSKIvEhrbt6hlOclb84vORW
AMiKvqSSJsaMufix+lZjOE5CmZRwVTvQFhKhagpfIWvjiVK3TGWGbDnoOFB9rQpIBRQAO6P+5trp
YY8L0tjQQ0tTelr8GTmc7ZGMchrlIYkF3xQ/2XfjE8wf1FzCWHVT3dz1bafgLe3yuIxxWCVBGbTS
lfU4aygEhYCi5o7t6NrZKn47qziuNFVFRryAFjRQNzoBlip2Y9dWDpBEwAV6CgZG/Nu9TizxRR1G
5Sjv3sv4v/OI0LyV5Sboytm0dandiMgJBMqSaI1fC7JCkzcYjPdC2GpdO0GuYmf6f2Kd+vIgZI8n
WSworkJdAr0xOJML4SOxEmrveL/k5TE9AAFPQywZ6aH7N7kt8aNY1+mQSkUo9nHKxMP60btx9YFr
4reCbP0Ju8M4bZc/5SZ5ncJXPZieTHXPS6TxUL3cN0j5N7acf9jomUhO8nHCnu0jFGvAdYZThDPf
5FNyQTR5kbvQTSSrORxT6KftC+Rhm709I/c1crfswIk9SuhIIf1bfTI9wU7/b3V4VcxO2k4MahZW
7CooPWxKzKc+eU9Pd2ATvwB9jymxDX/bzB5rm6nJPeNDtCUCZDk6n6jeq68fX+uHkjYFJLQmKo5B
rFLmDItI0FGoyw/vm5OycIuPX0BNh0dcW/A7sDL3cjsECj+KbZw4PGtLP2XDxULjU1ZYytqPZE8q
E+6nck9+v3izE5tZwnuaj4SIe5D2ucIfQmpQ4E+KX+vv7NgerY6hqx1ZEFAiJQzOqAOUISlvbS+b
mDvhLwI7af3p7I9cPkJ4izRsbPNI9zzAcj4x9mWAqzkniBVv9Jnhq1ps/r9OqVQhKbh+9fZVB6x7
QcZB3PJMmQlvSprbDqfQkXzzCPTrfoVw2mDCgllIACLfYxtL1cTLE2eoVkb1CTU1GbJ5SXr0XRAN
bIWRtc17eXWBZD4BDJFj42ESyyjgNJ2JT4gEiI/hl80A2rBYz3HK807FDm8shTL1qacsAmv3aN+k
mw4dYsg3H0QSgbF5N2q+pR0hM08tWpomDTMBp0bYWxo+RJJCKToTKUKkrGcCMvUccyNnzKAp6Jvo
rZO+8gPEPxV4mJShnjNIEYjiv1OryFydaEsUfF/FqT/pK3RUX37lvpXALaDFJm+t1/0s330xM1eh
aDZrQpt/psg5oqvN88nHiMgaDfvfIAY9I8tUDHVYAtgkiwRiDNE+ovHlTAJi3gKH3gKxZL7eQkZF
c1lgDYVU92TGRFFl3IHuL8OXcIP3bfNTZhTZ9beuWcZu6yHski3Um94upkcTBJ6F3OZE4yxpPSz6
CF0gRlPkuDClEx59f+F52WrKo6QALHPXbUT2Ujr7Bpvl9aCgYcnGZiDzMRnpaXX8FTx7mPyCmVuM
N1FpOOu7gY3dhEaKacFDB+1kjcpL/tkoT0fii98dIvyEvK1a7J3esFEnWLY6jiKJe7zU0iz8Wf/c
5OkM0sYuMcdcAGcZGNneiq+XiOPPsH2FZ74kxoaYtZm0Ch5HO/tQ0fJP1GsJFjmE5p9+goyCwh13
uu5C+sYj6jujxevZWUIco9lrDKJ/aQhkeHYPY34KxSoHTA9QuJFZg0LSNS3/bKp6nw7qsAONmn1Y
Q3gAPOhL8X3fD2p83WiBe/7H5d4GoDUGngpMU/4YVmpBo2XcfuQiq35x7EwKnj465VEocAVguAg8
7kq+d28WrhbpGDXp3qoWVwZBA1wVywH0X83/IXSkrjNYQQ+47dSsIZZ8httycZw8Md9tC1QxsRvA
IZ9PuGWsOpSKjLI1Fn1EGgiiKACJdgxjUndTNqikS7TXQbKVOYJ2ruZu4rDnr0JVq35D9D+f9gCN
PsdpAyp4Uyl1nwpGeryQUPIgHDuGANJhe5ZUlFlPFiMrW4wqxJ06JmqhIdhVlI71j6LOPYXH/bSi
PSSC4eDX9mawFku4WBYTm8faIBhfImbe7zkd9+Y3En2aucwpeOlc3MUeeLmP50vOrRS+Hqzlb4Fn
XFvg5K1/f5oZVOo6ure1yAqWmxIjM7irOjylqchgNm4i7eNdZNPXgJwtKiYNuHrhmiNk2WDMNngB
Ada+bS0R3GvOQYt/00qQMgqzTJVlnQpg8/nP5Aks1pUAnxjofGngx9h+ymv0ait6np6cHPpXEtKw
+ImAOx59qocrgsW3KyIxET6khcZ8oh3JzMvFFnBMkkxjatEd+8N0F+VNVc+XR3TnnsxsNr0N9Bds
dZi79Q6h150FPLRuA/tU9ZdTwTlfa7UIaC6UulN6DfsNFA3ISe1B+jAGeIGofhCTjQkvbcrwiY49
fa2HnEgsk5euznD63DClSVZ8MqwrTxeZycZN05R9WdvbjAcvU4BnVkDjMY8LhwQOQuVaIhvajs1q
fYzAJdcXRmKBBN+c6cID44mZ25srXka2OtkVjM1+torsuuGCGw+dTcwmsZ2+ONiiq6f957JYtmey
Ujb/F+0A8dYMlBoF2v5yJD8gCqPxpVMdyPi7KRgxiwoPOyHeZXX9hG/MeidhVV/XxC9cqIgyjK6x
P9CXooCp2p5Vw19qxddIuH4OpxPLUfRO/+9n8GGGwAE0IUqUb55dBTGJi728SZVXVwWP2Uwtu09v
MmZznSjV4XLlGR3TNWT0XAEoBCGFxiAgh9Ub2vn6tUTTnlbpZAFoL60hJlvNB+drlRmIvA12AlYt
bIpI0KzYw08sWKBgyP6hhTEyCJd1Adik8h0hOHtlTMaXEq+JfZun8kzoEHVvlCntaT9cPNXDM0+x
l83kk9jIT9PZUgiPo1nwQILPhW9R3sKOZo3ynIHNslkqH6JcCQk2ghZJ/TYZgij/BrdWxU1YWY0i
mA345FXVDNE8rgQSXWbmLXUGOVkmRPm4VAbQMg7sv0WwbPkzPFPWZInORGCf4hR/K5aZHcAQfxQc
eee84//aFfVP9swpD67gXXMQY/CUmfHMjAKmmYDZUDX63CVW5Ub/FXYRpm0ZNh39jK7nX/hbIg0z
80ophM6qXN8/u/GmU5N46oyC67XIY4ZutDWiPetjZF+Eiyg8KhDwfrWdNBwDhuIdAjGk76137XYq
+g3+aRz2nF7o7RaikjXAOGQWd0PymkWDp9hOb+B3bDkwNntsC0fYQAbSoIAwfs4VQ+qI0fXKsULu
MS81nyxqeQ36fOMYWsQ7fOf/+nnNbqkpUkgRN1ht31s3Yv19NKXhxubsZ0fBPbuniwiUpfd0i60+
xiOQlsoTXYnHA7nKhOH8QBaLAs5mLdxdEzTElgHh0ZM58vA/8IPQPPC+MXI/FytYbDlUgisXWa7X
zHRp0B1ze4ytNW3gKkp7H33nxMzVjPYsngcujaRb7H6bt7S/iY4R/mOwfypevchru+iCKDPs4N4j
hrbKpr72J+sR+1XB1rtVNyrRrg84YAw7bUkJrIMV9oviKQfXNaUK9CnqE5Hbp18fTubZYKnh7g+w
O8BfMo0wnBO3tl5JUZyuD2gVErznf1+dMf7NQ/J6oa+0MXR8pgE3Yx0zkmB0TcGbzjg615Fw8+Du
a1w/uHbE+xI73zDA1Ydz/ugseYH8otjMcfjMw825eZjjuOU7yS2bgUg3E30e5FXIoBGvcbaNaFQA
Ulb3dWHHCgaDp+AtZyuXysKUW/RpzmdC4tKo/4oiLjeuf3qk2eqVCpEHlrJDkFmRWSWwWQF8y8XL
H2yMqLcDyfZ5ngFp3qrPIpGK4zA02ZiAEmIXFagcD3WnhdbptTVh7wGSujbZGzk1Jyxf+GcSxPmz
R911K703VfGX8UFd4XhdqRVu7UYqa+SoddUwQX575RYa8vt1jrX+0TnX/yDXZFJV/0wT8O44QSCJ
S6W8k7aVf6Hjfo9IAKPHwvvCzH0HeE8n3ayRoUjb+oTM94rhAW+kwxZtZMNIy7FyupLnHdp50gzv
ubugGfeH7S3w59+/bK9v5Wnbzmcs9N0w9qYIOEnIWVSf4q+JYKbbSPB3A1EAkd/CYj368jcbOTNS
vf8U5S4sdZMP6ob3dpfTIaxwujmygaPTtsHdVEiwUym+GlHCl7gzurrlZ9Us8a8ft/6NZiQKMb2S
9U8yRMDiOFeaGdAdjs9W1zGDkCHLNXrRk9ouuc0IN/j7M6PjdGPvWlgy5/JKoAVKZIsThNGWHTPy
idITvvm0CAojeNH/xAey1fvR33uaxiGA4fLM4QO1Bag4ETbH/G0qXCtwU/qIqaB0vIbwMLsmKF8h
zAUKruyRmy/5bezQZK7+3IUzAkuLY3naGCtdMYiwkkDbHP9UavfR0Zce6+hPGPxebxQdw15pP/7W
AUHJkgUcZel7Q7GEL4P79mRwAP/P6FnfwpVLzz0vKZHfBsHuHyJL0uyhTKBtaeKsnQ/+UfezRyHb
llT/7cz4loEnx/Pi5mNz4H359NNNDIlxwfMk/RmRVlG+asb1zpQipBmdL0p9mtgzUgHIUClkmIfT
9JlZvufiKe/WvurIquqSPHslyoidXGtYKvfwc8ei+paYZIBkzzZfCQ+8JiytZiUpCCD3/D8LPyJk
9PV4ZWUzQeAOe+SG0824Q1ntWWoaF8z4nTdS/rPbTPkY7vfWYL5ONJ0mz4lc838sGTgoH0q2BRjl
Z7zCckAZabt7WTCup008QdIWpPGSFnhjgWRE5XvygrS0iKMyTPC5xJ4wWIyeVKcf46NJee5RB+yD
C9YDITQmVUXJbWCpDbU6ta+st3BsCCgYfXyuqnX1xBsryL5Ogslam+a7Q1QH6W4/Vu1qR8WyBfTy
gxAyezXRZfnuTyk/siTbKeegxhdLsDGf7PbWz6o6Bk2hPDP9/nMKDdacyMgB35YRlLS86/idTjsN
aL1lZtG6ZKL+2fPGmF5yMiNRZZRBN5HwUBumaFp81e/1Nm4PbVgFB/mbkT6tTm81m7Zwdlu8Bt/k
2F8pNcJcn6PXvyCvuVy3tHts98QTenMbDrJwGRM2otrgUjzZA2mD44DqcKPOYKUadRYtahBNX/PK
bP7FLyheWlyZsIZjKFk200mbNIvhNmYvUEwECh9GC2Ij/1o2cnHK8vLla33drXEDygP7pGLy7ZR3
J/FHVqEv5xmG6KCAv5yBVecEXd0VDBvVlrQx/n2mfrslELw67IBYQyXN+IUhw6On5+kfJBiSmEhi
FNvYSu4lABcYSMZkdyCKfIL/FqtXBGt25bXzlpOWAEKCvQmPQZigZpnk7HIgy/UUP8puEzarJDYV
n8N23asrqScmfFEWZcEWn9FOJCNxB0+zlMhUWuioxaCRoztm9EhV3JfEdtFGqViUjResuamZxufg
71/Gk0Yq/J33Byj/lDku35UaYd/oograUEE6NNAjpf8w94a7eXVGdAKT/rWpIfVXiQphgl+dhA4G
DQR5B3RibhiiBoONOOmULru2Ai0ly06DCRfzc5knOf2OoLUqFXxcWGBftmAc9EW86h9CcWLCe5Ix
HSF37kIqyWg8OcWBCrJIWAegI3BGSPt+t6jz17pXi0imEIlFbfQJQ4nhr62DEgrgLuBoJIT/PSyt
dzfMuJ/7c7J/JYMZ28Ibg4JELvAzeQRxHNZU7FQwP/erc1pfA2K2XZtVV/09e0WuAI807bVmevya
BCxkP+mnsW6FWMjRpTDiynivMFeH1jmUnVzGiqOaYfvowQ2/LKJeQKqhzeJjW3RPvBz+ortgrN8k
rzra60mPPQUbc16tTWipO2mMyPXk+iZhMulCp4NECDX3XMKOWDlzHZx7tIhJPWiGVzasK57Vg9nt
fLTSSZ+z2AarlNy6axvPj+eaUsn6VSzJZ12j7OYUfT3UUtot3J0ANMxaTDSYsAivmEbGgq/6jciK
kTMX+4IEUEkVRbgOrZQxZqFNS3acOTm9By2ong069+JHyTegly7F6krGl2xFgd20hA8TvSrCI1S9
a6VjZzU1+zjTushY5g/sSOvEK56bRZP50qNmhHdKzqU0/3YMdBP7M/drDkDvBNaEChjFsXMJc7T5
TbwLiZRfijk+KKv9M+hzCxGxyvFxw8akT5OTG04zIBW97/a4pNgLImGMnur2xfItet5jSBS7cyhK
zFSwiD6d8fKfMY6FG7G/GFT8nWdxMcV6RjeMixzrzTHGnErkbVZL0K4Bdn7YT9pY7Tn7/En4vHr3
v74lKiZ/y2nt8gT1zwcJr/NO+6FfIlgHLV9dZ5/XRaEwsoQcCbomRamJMhcr+wDoouwLNMHl6AWt
u9TXag/qJMoAO2xjZ0R3SnIhprLNv5QfaFZcYh/0wQuNsH1JBP9KqKbP4HzCG9FllBVDHbinHmmZ
8cpkWA==
`pragma protect end_protected
